module interconect_cells(
	clk,
	reset,
	divisor,
	dividend,
	mode,
	valid_input,
	valid_output,
	final_output
);

	input [31:0] dividend;
	input [15:0] divisor;

	input clk, reset;
	input valid_input, mode;

	output valid_output;
	output [17:0] final_output;

	reg [16:0] div_res;
	reg [15:0] mod_res;

	wire [16:0] wire_out_quotient;
	wire [14:0] wire_out_remainder;

	wire one=1'b1;

	always @(*) begin
		if (reset) begin
			div_res[16] = 'd0;
			div_res[15] = 'd0;
			div_res[14] = 'd0;
			div_res[13] = 'd0;
			div_res[12] = 'd0;
			div_res[11] = 'd0;
			div_res[10] = 'd0;
			div_res[9] = 'd0;
			div_res[8] = 'd0;
			div_res[7] = 'd0;
			div_res[6] = 'd0;
			div_res[5] = 'd0;
			div_res[4] = 'd0;
			div_res[3] = 'd0;
			div_res[2] = 'd0;
			div_res[1] = 'd0;
			div_res[0] = 'd0;
		end else begin
			div_res[16] = ~wire_out_quotient[16];
			div_res[15] = ~wire_out_quotient[15];
			div_res[14] = ~wire_out_quotient[14];
			div_res[13] = ~wire_out_quotient[13];
			div_res[12] = ~wire_out_quotient[12];
			div_res[11] = ~wire_out_quotient[11];
			div_res[10] = ~wire_out_quotient[10];
			div_res[9] = ~wire_out_quotient[9];
			div_res[8] = ~wire_out_quotient[8];
			div_res[7] = ~wire_out_quotient[7];
			div_res[6] = ~wire_out_quotient[6];
			div_res[5] = ~wire_out_quotient[5];
			div_res[4] = ~wire_out_quotient[4];
			div_res[3] = ~wire_out_quotient[3];
			div_res[2] = ~wire_out_quotient[2];
			div_res[1] = ~wire_out_quotient[1];
			div_res[0] = ~wire_out_quotient[0];
		end
	end

	always @(*) begin
		if (reset) begin
			mod_res[15] ='d0;
			mod_res[14] ='d0;
			mod_res[13] ='d0;
			mod_res[12] ='d0;
			mod_res[11] ='d0;
			mod_res[10] ='d0;
			mod_res[9] = 'd0;
			mod_res[8] = 'd0;
			mod_res[7] = 'd0;
			mod_res[6] = 'd0;
			mod_res[5] = 'd0;
			mod_res[4] = 'd0;
			mod_res[3] = 'd0;
			mod_res[2] = 'd0;
			mod_res[1] = 'd0;
			mod_res[0] = 'd0;	
		end else begin
			mod_res[15] = wire_out_quotient[0];
			mod_res[14] = wire_out_remainder[14];
			mod_res[13] = wire_out_remainder[13];
			mod_res[12] = wire_out_remainder[12];
			mod_res[11] = wire_out_remainder[11];
			mod_res[10] = wire_out_remainder[10];
			mod_res[9] = wire_out_remainder[9];
			mod_res[8] = wire_out_remainder[8];
			mod_res[7] = wire_out_remainder[7];
			mod_res[6] = wire_out_remainder[6];
			mod_res[5] = wire_out_remainder[5];
			mod_res[4] = wire_out_remainder[4];
			mod_res[3] = wire_out_remainder[3];
			mod_res[2] = wire_out_remainder[2];
			mod_res[1] = wire_out_remainder[1];
			mod_res[0] = wire_out_remainder[0];	
		end
	end

	always @(*) begin
		if (mod_res[15] == 1) begin
			mod_res = mod_res + divisor;
		end
	end

	assign final_output = (mode) ? div_res : mod_res;

	//div_cell cas_X_Y (T_in,Divisor_in,Remainder_in/dividend,Remainder_out,C_in,C_out);
	//1st row
	div_cell cas_0_15 ( one ,  divisor[15] ,  dividend[31] ,   wire_out_quotient[16] ,  wire_0_14_15_curry ,  hang_0_wire_15 );

	div_cell cas_0_14 ( one ,  divisor[14] ,  dividend[30] ,  wire_0_14_1_15_remainter ,  wire_0_13_14_curry ,  wire_0_14_15_curry );
	div_cell cas_0_13 ( one ,  divisor[13] ,  dividend[29] ,  wire_0_13_1_14_remainter ,  wire_0_12_13_curry ,  wire_0_13_14_curry );
	div_cell cas_0_12 ( one ,  divisor[12] ,  dividend[28] ,  wire_0_12_1_13_remainter ,  wire_0_11_12_curry ,  wire_0_12_13_curry );
	div_cell cas_0_11 ( one ,  divisor[11] ,  dividend[27] ,  wire_0_11_1_12_remainter ,  wire_0_10_11_curry ,  wire_0_11_12_curry );
	div_cell cas_0_10 ( one ,  divisor[10] ,  dividend[26] ,  wire_0_10_1_11_remainter ,  wire_0_09_10_curry ,  wire_0_10_11_curry );
	div_cell cas_0_9 ( one ,  divisor[9] ,  dividend[25] ,  wire_0_9_1_10_remainter ,  wire_0_08_09_curry ,  wire_0_09_10_curry );
	div_cell cas_0_8 ( one ,  divisor[8] ,  dividend[24] ,  wire_0_8_1_9_remainter ,  wire_0_07_08_curry ,  wire_0_08_09_curry );
	div_cell cas_0_7 ( one ,  divisor[7] ,  dividend[23] ,  wire_0_7_1_8_remainter ,  wire_0_06_07_curry ,  wire_0_07_08_curry );
	div_cell cas_0_6 ( one ,  divisor[6] ,  dividend[22] ,  wire_0_6_1_7_remainter ,  wire_0_05_06_curry ,  wire_0_06_07_curry );
	div_cell cas_0_5 ( one ,  divisor[5] ,  dividend[21] ,  wire_0_5_1_6_remainter ,  wire_0_04_05_curry ,  wire_0_05_06_curry );
	div_cell cas_0_4 ( one ,  divisor[4] ,  dividend[20] ,  wire_0_4_1_5_remainter ,  wire_0_03_04_curry ,  wire_0_04_05_curry );
	div_cell cas_0_3 ( one ,  divisor[3] ,  dividend[19] ,  wire_0_3_1_4_remainter ,  wire_0_02_03_curry ,  wire_0_03_04_curry );
	div_cell cas_0_2 ( one ,  divisor[2] ,  dividend[18] ,  wire_0_2_1_3_remainter ,  wire_0_01_02_curry ,  wire_0_02_03_curry );
	div_cell cas_0_1 ( one ,  divisor[1] ,  dividend[17] ,  wire_0_1_1_2_remainter ,  wire_0_00_01_curry ,  wire_0_01_02_curry );

	div_cell cas_0_0 ( one ,  divisor[0] ,  dividend[16] ,  wire_0_0_1_1_remainter ,  one ,  wire_0_00_01_curry );

	//div_cell cas_X_Y (T_in,Divisor_in,Remainder_in/dividend,Remainder_out,C_in,C_out);
	//2nd row
	div_cell cas_1_15 (~wire_out_quotient[16], divisor[15], wire_0_14_1_15_remainter,  wire_out_quotient[15], wire_1_14_15_curry, hang_1_wire_15);

	div_cell cas_1_14 ( ~wire_out_quotient[16] ,  divisor[14] ,  wire_0_13_1_14_remainter ,  wire_1_14_2_15_remainter ,  wire_1_13_14_curry ,  wire_1_14_15_curry );
	div_cell cas_1_13 ( ~wire_out_quotient[16] ,  divisor[13] ,  wire_0_12_1_13_remainter ,  wire_1_13_2_14_remainter ,  wire_1_12_13_curry ,  wire_1_13_14_curry );
	div_cell cas_1_12 ( ~wire_out_quotient[16] ,  divisor[12] ,  wire_0_11_1_12_remainter ,  wire_1_12_2_13_remainter ,  wire_1_11_12_curry ,  wire_1_12_13_curry );
	div_cell cas_1_11 ( ~wire_out_quotient[16] ,  divisor[11] ,  wire_0_10_1_11_remainter ,  wire_1_11_2_12_remainter ,  wire_1_10_11_curry ,  wire_1_11_12_curry );
	div_cell cas_1_10 ( ~wire_out_quotient[16] ,  divisor[10] ,  wire_0_9_1_10_remainter ,  wire_1_10_2_11_remainter ,  wire_1_09_10_curry ,  wire_1_10_11_curry );
	div_cell cas_1_9 ( ~wire_out_quotient[16] ,  divisor[9] ,  wire_0_8_1_9_remainter ,  wire_1_9_2_10_remainter ,  wire_1_08_09_curry ,  wire_1_09_10_curry );
	div_cell cas_1_8 ( ~wire_out_quotient[16] ,  divisor[8] ,  wire_0_7_1_8_remainter ,  wire_1_8_2_9_remainter ,  wire_1_07_08_curry ,  wire_1_08_09_curry );
	div_cell cas_1_7 ( ~wire_out_quotient[16] ,  divisor[7] ,  wire_0_6_1_7_remainter ,  wire_1_7_2_8_remainter ,  wire_1_06_07_curry ,  wire_1_07_08_curry );
	div_cell cas_1_6 ( ~wire_out_quotient[16] ,  divisor[6] ,  wire_0_5_1_6_remainter ,  wire_1_6_2_7_remainter ,  wire_1_05_06_curry ,  wire_1_06_07_curry );
	div_cell cas_1_5 ( ~wire_out_quotient[16] ,  divisor[5] ,  wire_0_4_1_5_remainter ,  wire_1_5_2_6_remainter ,  wire_1_04_05_curry ,  wire_1_05_06_curry );
	div_cell cas_1_4 ( ~wire_out_quotient[16] ,  divisor[4] ,  wire_0_3_1_4_remainter ,  wire_1_4_2_5_remainter ,  wire_1_03_04_curry ,  wire_1_04_05_curry );
	div_cell cas_1_3 ( ~wire_out_quotient[16] ,  divisor[3] ,  wire_0_2_1_3_remainter ,  wire_1_3_2_4_remainter ,  wire_1_02_03_curry ,  wire_1_03_04_curry );
	div_cell cas_1_2 ( ~wire_out_quotient[16] ,  divisor[2] ,  wire_0_1_1_2_remainter ,  wire_1_2_2_3_remainter ,  wire_1_01_02_curry ,  wire_1_02_03_curry );
	div_cell cas_1_1 ( ~wire_out_quotient[16] ,  divisor[1] ,  wire_0_0_1_1_remainter ,  wire_1_1_2_2_remainter ,  wire_1_00_01_curry ,  wire_1_01_02_curry );

	div_cell cas_1_0 ( ~wire_out_quotient[16] ,  divisor[0] ,  dividend[15] ,  wire_1_0_2_1_remainter ,  ~wire_out_quotient[16] ,  wire_1_00_01_curry );

	//3rd row
	div_cell cas_2_15 ( ~wire_out_quotient[15] ,  divisor[15] ,  wire_1_14_2_15_remainter ,   wire_out_quotient[14] ,  wire_2_14_15_curry ,  hang_2_wire_15 );

	div_cell cas_2_14 ( ~wire_out_quotient[15] ,  divisor[14] ,  wire_1_13_2_14_remainter ,  wire_2_14_3_15_remainter ,  wire_2_13_14_curry ,  wire_2_14_15_curry );
	div_cell cas_2_13 ( ~wire_out_quotient[15] ,  divisor[13] ,  wire_1_12_2_13_remainter ,  wire_2_13_3_14_remainter ,  wire_2_12_13_curry ,  wire_2_13_14_curry );
	div_cell cas_2_12 ( ~wire_out_quotient[15] ,  divisor[12] ,  wire_1_11_2_12_remainter ,  wire_2_12_3_13_remainter ,  wire_2_11_12_curry ,  wire_2_12_13_curry );
	div_cell cas_2_11 ( ~wire_out_quotient[15] ,  divisor[11] ,  wire_1_10_2_11_remainter ,  wire_2_11_3_12_remainter ,  wire_2_10_11_curry ,  wire_2_11_12_curry );
	div_cell cas_2_10 ( ~wire_out_quotient[15] ,  divisor[10] ,  wire_1_9_2_10_remainter ,  wire_2_10_3_11_remainter ,  wire_2_09_10_curry ,  wire_2_10_11_curry );
	div_cell cas_2_9 ( ~wire_out_quotient[15] ,  divisor[9] ,  wire_1_8_2_9_remainter ,  wire_2_9_3_10_remainter ,  wire_2_08_09_curry ,  wire_2_09_10_curry );
	div_cell cas_2_8 ( ~wire_out_quotient[15] ,  divisor[8] ,  wire_1_7_2_8_remainter ,  wire_2_8_3_9_remainter ,  wire_2_07_08_curry ,  wire_2_08_09_curry );
	div_cell cas_2_7 ( ~wire_out_quotient[15] ,  divisor[7] ,  wire_1_6_2_7_remainter ,  wire_2_7_3_8_remainter ,  wire_2_06_07_curry ,  wire_2_07_08_curry );
	div_cell cas_2_6 ( ~wire_out_quotient[15] ,  divisor[6] ,  wire_1_5_2_6_remainter ,  wire_2_6_3_7_remainter ,  wire_2_05_06_curry ,  wire_2_06_07_curry );
	div_cell cas_2_5 ( ~wire_out_quotient[15] ,  divisor[5] ,  wire_1_4_2_5_remainter ,  wire_2_5_3_6_remainter ,  wire_2_04_05_curry ,  wire_2_05_06_curry );
	div_cell cas_2_4 ( ~wire_out_quotient[15] ,  divisor[4] ,  wire_1_3_2_4_remainter ,  wire_2_4_3_5_remainter ,  wire_2_03_04_curry ,  wire_2_04_05_curry );
	div_cell cas_2_3 ( ~wire_out_quotient[15] ,  divisor[3] ,  wire_1_2_2_3_remainter ,  wire_2_3_3_4_remainter ,  wire_2_02_03_curry ,  wire_2_03_04_curry );
	div_cell cas_2_2 ( ~wire_out_quotient[15] ,  divisor[2] ,  wire_1_1_2_2_remainter ,  wire_2_2_3_3_remainter ,  wire_2_01_02_curry ,  wire_2_02_03_curry );
	div_cell cas_2_1 ( ~wire_out_quotient[15] ,  divisor[1] ,  wire_1_0_2_1_remainter ,  wire_2_1_3_2_remainter ,  wire_2_00_01_curry ,  wire_2_01_02_curry );

	div_cell cas_2_0 ( ~wire_out_quotient[15] ,  divisor[0] ,  dividend[14] ,  wire_2_0_3_1_remainter ,  ~wire_out_quotient[15] ,  wire_2_00_01_curry );

	//4th row
	div_cell cas_3_15 ( ~wire_out_quotient[14] ,  divisor[15] ,  wire_2_14_3_15_remainter ,   wire_out_quotient[13] ,  wire_3_14_15_curry ,  hang_3_wire_15 );

	div_cell cas_3_14 ( ~wire_out_quotient[14] ,  divisor[14] ,  wire_2_13_3_14_remainter ,  wire_3_14_4_15_remainter ,  wire_3_13_14_curry ,  wire_3_14_15_curry );
	div_cell cas_3_13 ( ~wire_out_quotient[14] ,  divisor[13] ,  wire_2_12_3_13_remainter ,  wire_3_13_4_14_remainter ,  wire_3_12_13_curry ,  wire_3_13_14_curry );
	div_cell cas_3_12 ( ~wire_out_quotient[14] ,  divisor[12] ,  wire_2_11_3_12_remainter ,  wire_3_12_4_13_remainter ,  wire_3_11_12_curry ,  wire_3_12_13_curry );
	div_cell cas_3_11 ( ~wire_out_quotient[14] ,  divisor[11] ,  wire_2_10_3_11_remainter ,  wire_3_11_4_12_remainter ,  wire_3_10_11_curry ,  wire_3_11_12_curry );
	div_cell cas_3_10 ( ~wire_out_quotient[14] ,  divisor[10] ,  wire_2_9_3_10_remainter ,  wire_3_10_4_11_remainter ,  wire_3_09_10_curry ,  wire_3_10_11_curry );
	div_cell cas_3_9 ( ~wire_out_quotient[14] ,  divisor[9] ,  wire_2_8_3_9_remainter ,  wire_3_9_4_10_remainter ,  wire_3_08_09_curry ,  wire_3_09_10_curry );
	div_cell cas_3_8 ( ~wire_out_quotient[14] ,  divisor[8] ,  wire_2_7_3_8_remainter ,  wire_3_8_4_9_remainter ,  wire_3_07_08_curry ,  wire_3_08_09_curry );
	div_cell cas_3_7 ( ~wire_out_quotient[14] ,  divisor[7] ,  wire_2_6_3_7_remainter ,  wire_3_7_4_8_remainter ,  wire_3_06_07_curry ,  wire_3_07_08_curry );
	div_cell cas_3_6 ( ~wire_out_quotient[14] ,  divisor[6] ,  wire_2_5_3_6_remainter ,  wire_3_6_4_7_remainter ,  wire_3_05_06_curry ,  wire_3_06_07_curry );
	div_cell cas_3_5 ( ~wire_out_quotient[14] ,  divisor[5] ,  wire_2_4_3_5_remainter ,  wire_3_5_4_6_remainter ,  wire_3_04_05_curry ,  wire_3_05_06_curry );
	div_cell cas_3_4 ( ~wire_out_quotient[14] ,  divisor[4] ,  wire_2_3_3_4_remainter ,  wire_3_4_4_5_remainter ,  wire_3_03_04_curry ,  wire_3_04_05_curry );
	div_cell cas_3_3 ( ~wire_out_quotient[14] ,  divisor[3] ,  wire_2_2_3_3_remainter ,  wire_3_3_4_4_remainter ,  wire_3_02_03_curry ,  wire_3_03_04_curry );
	div_cell cas_3_2 ( ~wire_out_quotient[14] ,  divisor[2] ,  wire_2_1_3_2_remainter ,  wire_3_2_4_3_remainter ,  wire_3_01_02_curry ,  wire_3_02_03_curry );
	div_cell cas_3_1 ( ~wire_out_quotient[14] ,  divisor[1] ,  wire_2_0_3_1_remainter ,  wire_3_1_4_2_remainter ,  wire_3_00_01_curry ,  wire_3_01_02_curry );

	div_cell cas_3_0 ( ~wire_out_quotient[14] ,  divisor[0] ,  dividend[13] ,  wire_3_0_4_1_remainter ,  ~wire_out_quotient[14] ,  wire_3_00_01_curry );

	//5th row
	div_cell cas_4_15 ( ~wire_out_quotient[13] ,  divisor[15] ,  wire_3_14_4_15_remainter ,   wire_out_quotient[12] ,  wire_4_14_15_curry ,  hang_4_wire_15 );

	div_cell cas_4_14 ( ~wire_out_quotient[13] ,  divisor[14] ,  wire_3_13_4_14_remainter ,  wire_4_14_5_15_remainter ,  wire_4_13_14_curry ,  wire_4_14_15_curry );
	div_cell cas_4_13 ( ~wire_out_quotient[13] ,  divisor[13] ,  wire_3_12_4_13_remainter ,  wire_4_13_5_14_remainter ,  wire_4_12_13_curry ,  wire_4_13_14_curry );
	div_cell cas_4_12 ( ~wire_out_quotient[13] ,  divisor[12] ,  wire_3_11_4_12_remainter ,  wire_4_12_5_13_remainter ,  wire_4_11_12_curry ,  wire_4_12_13_curry );
	div_cell cas_4_11 ( ~wire_out_quotient[13] ,  divisor[11] ,  wire_3_10_4_11_remainter ,  wire_4_11_5_12_remainter ,  wire_4_10_11_curry ,  wire_4_11_12_curry );
	div_cell cas_4_10 ( ~wire_out_quotient[13] ,  divisor[10] ,  wire_3_9_4_10_remainter ,  wire_4_10_5_11_remainter ,  wire_4_09_10_curry ,  wire_4_10_11_curry );
	div_cell cas_4_9 ( ~wire_out_quotient[13] ,  divisor[9] ,  wire_3_8_4_9_remainter ,  wire_4_9_5_10_remainter ,  wire_4_08_09_curry ,  wire_4_09_10_curry );
	div_cell cas_4_8 ( ~wire_out_quotient[13] ,  divisor[8] ,  wire_3_7_4_8_remainter ,  wire_4_8_5_9_remainter ,  wire_4_07_08_curry ,  wire_4_08_09_curry );
	div_cell cas_4_7 ( ~wire_out_quotient[13] ,  divisor[7] ,  wire_3_6_4_7_remainter ,  wire_4_7_5_8_remainter ,  wire_4_06_07_curry ,  wire_4_07_08_curry );
	div_cell cas_4_6 ( ~wire_out_quotient[13] ,  divisor[6] ,  wire_3_5_4_6_remainter ,  wire_4_6_5_7_remainter ,  wire_4_05_06_curry ,  wire_4_06_07_curry );
	div_cell cas_4_5 ( ~wire_out_quotient[13] ,  divisor[5] ,  wire_3_4_4_5_remainter ,  wire_4_5_5_6_remainter ,  wire_4_04_05_curry ,  wire_4_05_06_curry );
	div_cell cas_4_4 ( ~wire_out_quotient[13] ,  divisor[4] ,  wire_3_3_4_4_remainter ,  wire_4_4_5_5_remainter ,  wire_4_03_04_curry ,  wire_4_04_05_curry );
	div_cell cas_4_3 ( ~wire_out_quotient[13] ,  divisor[3] ,  wire_3_2_4_3_remainter ,  wire_4_3_5_4_remainter ,  wire_4_02_03_curry ,  wire_4_03_04_curry );
	div_cell cas_4_2 ( ~wire_out_quotient[13] ,  divisor[2] ,  wire_3_1_4_2_remainter ,  wire_4_2_5_3_remainter ,  wire_4_01_02_curry ,  wire_4_02_03_curry );
	div_cell cas_4_1 ( ~wire_out_quotient[13] ,  divisor[1] ,  wire_3_0_4_1_remainter ,  wire_4_1_5_2_remainter ,  wire_4_00_01_curry ,  wire_4_01_02_curry );

	div_cell cas_4_0 ( ~wire_out_quotient[13] ,  divisor[0] ,  dividend[12] ,  wire_4_0_5_1_remainter ,  ~wire_out_quotient[13] ,  wire_4_00_01_curry );

	//6th row
	div_cell cas_5_15 ( ~wire_out_quotient[12] ,  divisor[15] ,  wire_4_14_5_15_remainter ,   wire_out_quotient[11] ,  wire_5_14_15_curry ,  hang_5_wire_15 );

	div_cell cas_5_14 ( ~wire_out_quotient[12] ,  divisor[14] ,  wire_4_13_5_14_remainter ,  wire_5_14_6_15_remainter ,  wire_5_13_14_curry ,  wire_5_14_15_curry );
	div_cell cas_5_13 ( ~wire_out_quotient[12] ,  divisor[13] ,  wire_4_12_5_13_remainter ,  wire_5_13_6_14_remainter ,  wire_5_12_13_curry ,  wire_5_13_14_curry );
	div_cell cas_5_12 ( ~wire_out_quotient[12] ,  divisor[12] ,  wire_4_11_5_12_remainter ,  wire_5_12_6_13_remainter ,  wire_5_11_12_curry ,  wire_5_12_13_curry );
	div_cell cas_5_11 ( ~wire_out_quotient[12] ,  divisor[11] ,  wire_4_10_5_11_remainter ,  wire_5_11_6_12_remainter ,  wire_5_10_11_curry ,  wire_5_11_12_curry );
	div_cell cas_5_10 ( ~wire_out_quotient[12] ,  divisor[10] ,  wire_4_9_5_10_remainter ,  wire_5_10_6_11_remainter ,  wire_5_09_10_curry ,  wire_5_10_11_curry );
	div_cell cas_5_9 ( ~wire_out_quotient[12] ,  divisor[9] ,  wire_4_8_5_9_remainter ,  wire_5_9_6_10_remainter ,  wire_5_08_09_curry ,  wire_5_09_10_curry );
	div_cell cas_5_8 ( ~wire_out_quotient[12] ,  divisor[8] ,  wire_4_7_5_8_remainter ,  wire_5_8_6_9_remainter ,  wire_5_07_08_curry ,  wire_5_08_09_curry );
	div_cell cas_5_7 ( ~wire_out_quotient[12] ,  divisor[7] ,  wire_4_6_5_7_remainter ,  wire_5_7_6_8_remainter ,  wire_5_06_07_curry ,  wire_5_07_08_curry );
	div_cell cas_5_6 ( ~wire_out_quotient[12] ,  divisor[6] ,  wire_4_5_5_6_remainter ,  wire_5_6_6_7_remainter ,  wire_5_05_06_curry ,  wire_5_06_07_curry );
	div_cell cas_5_5 ( ~wire_out_quotient[12] ,  divisor[5] ,  wire_4_4_5_5_remainter ,  wire_5_5_6_6_remainter ,  wire_5_04_05_curry ,  wire_5_05_06_curry );
	div_cell cas_5_4 ( ~wire_out_quotient[12] ,  divisor[4] ,  wire_4_3_5_4_remainter ,  wire_5_4_6_5_remainter ,  wire_5_03_04_curry ,  wire_5_04_05_curry );
	div_cell cas_5_3 ( ~wire_out_quotient[12] ,  divisor[3] ,  wire_4_2_5_3_remainter ,  wire_5_3_6_4_remainter ,  wire_5_02_03_curry ,  wire_5_03_04_curry );
	div_cell cas_5_2 ( ~wire_out_quotient[12] ,  divisor[2] ,  wire_4_1_5_2_remainter ,  wire_5_2_6_3_remainter ,  wire_5_01_02_curry ,  wire_5_02_03_curry );
	div_cell cas_5_1 ( ~wire_out_quotient[12] ,  divisor[1] ,  wire_4_0_5_1_remainter ,  wire_5_1_6_2_remainter ,  wire_5_00_01_curry ,  wire_5_01_02_curry );

	div_cell cas_5_0 ( ~wire_out_quotient[12] ,  divisor[0] ,  dividend[11] ,  wire_5_0_6_1_remainter ,  ~wire_out_quotient[12] ,  wire_5_00_01_curry );

	//7th row
	div_cell cas_6_15 ( ~wire_out_quotient[11] ,  divisor[15] ,  wire_5_14_6_15_remainter ,   wire_out_quotient[10] ,  wire_6_14_15_curry ,  hang_6_wire_15 );

	div_cell cas_6_14 ( ~wire_out_quotient[11] ,  divisor[14] ,  wire_5_13_6_14_remainter ,  wire_6_14_7_15_remainter ,  wire_6_13_14_curry ,  wire_6_14_15_curry );
	div_cell cas_6_13 ( ~wire_out_quotient[11] ,  divisor[13] ,  wire_5_12_6_13_remainter ,  wire_6_13_7_14_remainter ,  wire_6_12_13_curry ,  wire_6_13_14_curry );
	div_cell cas_6_12 ( ~wire_out_quotient[11] ,  divisor[12] ,  wire_5_11_6_12_remainter ,  wire_6_12_7_13_remainter ,  wire_6_11_12_curry ,  wire_6_12_13_curry );
	div_cell cas_6_11 ( ~wire_out_quotient[11] ,  divisor[11] ,  wire_5_10_6_11_remainter ,  wire_6_11_7_12_remainter ,  wire_6_10_11_curry ,  wire_6_11_12_curry );
	div_cell cas_6_10 ( ~wire_out_quotient[11] ,  divisor[10] ,  wire_5_9_6_10_remainter ,  wire_6_10_7_11_remainter ,  wire_6_09_10_curry ,  wire_6_10_11_curry );
	div_cell cas_6_9 ( ~wire_out_quotient[11] ,  divisor[9] ,  wire_5_8_6_9_remainter ,  wire_6_9_7_10_remainter ,  wire_6_08_09_curry ,  wire_6_09_10_curry );
	div_cell cas_6_8 ( ~wire_out_quotient[11] ,  divisor[8] ,  wire_5_7_6_8_remainter ,  wire_6_8_7_9_remainter ,  wire_6_07_08_curry ,  wire_6_08_09_curry );
	div_cell cas_6_7 ( ~wire_out_quotient[11] ,  divisor[7] ,  wire_5_6_6_7_remainter ,  wire_6_7_7_8_remainter ,  wire_6_06_07_curry ,  wire_6_07_08_curry );
	div_cell cas_6_6 ( ~wire_out_quotient[11] ,  divisor[6] ,  wire_5_5_6_6_remainter ,  wire_6_6_7_7_remainter ,  wire_6_05_06_curry ,  wire_6_06_07_curry );
	div_cell cas_6_5 ( ~wire_out_quotient[11] ,  divisor[5] ,  wire_5_4_6_5_remainter ,  wire_6_5_7_6_remainter ,  wire_6_04_05_curry ,  wire_6_05_06_curry );
	div_cell cas_6_4 ( ~wire_out_quotient[11] ,  divisor[4] ,  wire_5_3_6_4_remainter ,  wire_6_4_7_5_remainter ,  wire_6_03_04_curry ,  wire_6_04_05_curry );
	div_cell cas_6_3 ( ~wire_out_quotient[11] ,  divisor[3] ,  wire_5_2_6_3_remainter ,  wire_6_3_7_4_remainter ,  wire_6_02_03_curry ,  wire_6_03_04_curry );
	div_cell cas_6_2 ( ~wire_out_quotient[11] ,  divisor[2] ,  wire_5_1_6_2_remainter ,  wire_6_2_7_3_remainter ,  wire_6_01_02_curry ,  wire_6_02_03_curry );
	div_cell cas_6_1 ( ~wire_out_quotient[11] ,  divisor[1] ,  wire_5_0_6_1_remainter ,  wire_6_1_7_2_remainter ,  wire_6_00_01_curry ,  wire_6_01_02_curry );

	div_cell cas_6_0 ( ~wire_out_quotient[11] ,  divisor[0] ,  dividend[10] ,  wire_6_0_7_1_remainter ,  ~wire_out_quotient[11] ,  wire_6_00_01_curry );

	//8th row
	div_cell cas_7_15 ( ~wire_out_quotient[10] ,  divisor[15] ,  wire_6_14_7_15_remainter ,   wire_out_quotient[9] ,  wire_7_14_15_curry ,  hang_7_wire_15 );

	div_cell cas_7_14 ( ~wire_out_quotient[10] ,  divisor[14] ,  wire_6_13_7_14_remainter ,  wire_7_14_8_15_remainter ,  wire_7_13_14_curry ,  wire_7_14_15_curry );
	div_cell cas_7_13 ( ~wire_out_quotient[10] ,  divisor[13] ,  wire_6_12_7_13_remainter ,  wire_7_13_8_14_remainter ,  wire_7_12_13_curry ,  wire_7_13_14_curry );
	div_cell cas_7_12 ( ~wire_out_quotient[10] ,  divisor[12] ,  wire_6_11_7_12_remainter ,  wire_7_12_8_13_remainter ,  wire_7_11_12_curry ,  wire_7_12_13_curry );
	div_cell cas_7_11 ( ~wire_out_quotient[10] ,  divisor[11] ,  wire_6_10_7_11_remainter ,  wire_7_11_8_12_remainter ,  wire_7_10_11_curry ,  wire_7_11_12_curry );
	div_cell cas_7_10 ( ~wire_out_quotient[10] ,  divisor[10] ,  wire_6_9_7_10_remainter ,  wire_7_10_8_11_remainter ,  wire_7_09_10_curry ,  wire_7_10_11_curry );
	div_cell cas_7_9 ( ~wire_out_quotient[10] ,  divisor[9] ,  wire_6_8_7_9_remainter ,  wire_7_9_8_10_remainter ,  wire_7_08_09_curry ,  wire_7_09_10_curry );
	div_cell cas_7_8 ( ~wire_out_quotient[10] ,  divisor[8] ,  wire_6_7_7_8_remainter ,  wire_7_8_8_9_remainter ,  wire_7_07_08_curry ,  wire_7_08_09_curry );
	div_cell cas_7_7 ( ~wire_out_quotient[10] ,  divisor[7] ,  wire_6_6_7_7_remainter ,  wire_7_7_8_8_remainter ,  wire_7_06_07_curry ,  wire_7_07_08_curry );
	div_cell cas_7_6 ( ~wire_out_quotient[10] ,  divisor[6] ,  wire_6_5_7_6_remainter ,  wire_7_6_8_7_remainter ,  wire_7_05_06_curry ,  wire_7_06_07_curry );
	div_cell cas_7_5 ( ~wire_out_quotient[10] ,  divisor[5] ,  wire_6_4_7_5_remainter ,  wire_7_5_8_6_remainter ,  wire_7_04_05_curry ,  wire_7_05_06_curry );
	div_cell cas_7_4 ( ~wire_out_quotient[10] ,  divisor[4] ,  wire_6_3_7_4_remainter ,  wire_7_4_8_5_remainter ,  wire_7_03_04_curry ,  wire_7_04_05_curry );
	div_cell cas_7_3 ( ~wire_out_quotient[10] ,  divisor[3] ,  wire_6_2_7_3_remainter ,  wire_7_3_8_4_remainter ,  wire_7_02_03_curry ,  wire_7_03_04_curry );
	div_cell cas_7_2 ( ~wire_out_quotient[10] ,  divisor[2] ,  wire_6_1_7_2_remainter ,  wire_7_2_8_3_remainter ,  wire_7_01_02_curry ,  wire_7_02_03_curry );
	div_cell cas_7_1 ( ~wire_out_quotient[10] ,  divisor[1] ,  wire_6_0_7_1_remainter ,  wire_7_1_8_2_remainter ,  wire_7_00_01_curry ,  wire_7_01_02_curry );
	
	div_cell cas_7_0 ( ~wire_out_quotient[10] ,  divisor[0] ,  dividend[9] ,  wire_7_0_8_1_remainter ,  ~wire_out_quotient[10] ,  wire_7_00_01_curry );

	//9th row
	div_cell cas_8_15 ( ~wire_out_quotient[9] ,  divisor[15] ,  wire_7_14_8_15_remainter ,   wire_out_quotient[8] ,  wire_8_14_15_curry ,  hang_8_wire_15 );

	div_cell cas_8_14 ( ~wire_out_quotient[9] ,  divisor[14] ,  wire_7_13_8_14_remainter ,  wire_8_14_9_15_remainter ,  wire_8_13_14_curry ,  wire_8_14_15_curry );
	div_cell cas_8_13 ( ~wire_out_quotient[9] ,  divisor[13] ,  wire_7_12_8_13_remainter ,  wire_8_13_9_14_remainter ,  wire_8_12_13_curry ,  wire_8_13_14_curry );
	div_cell cas_8_12 ( ~wire_out_quotient[9] ,  divisor[12] ,  wire_7_11_8_12_remainter ,  wire_8_12_9_13_remainter ,  wire_8_11_12_curry ,  wire_8_12_13_curry );
	div_cell cas_8_11 ( ~wire_out_quotient[9] ,  divisor[11] ,  wire_7_10_8_11_remainter ,  wire_8_11_9_12_remainter ,  wire_8_10_11_curry ,  wire_8_11_12_curry );
	div_cell cas_8_10 ( ~wire_out_quotient[9] ,  divisor[10] ,  wire_7_9_8_10_remainter ,  wire_8_10_9_11_remainter ,  wire_8_09_10_curry ,  wire_8_10_11_curry );
	div_cell cas_8_9 ( ~wire_out_quotient[9] ,  divisor[9] ,  wire_7_8_8_9_remainter ,  wire_8_9_9_10_remainter ,  wire_8_08_09_curry ,  wire_8_09_10_curry );
	div_cell cas_8_8 ( ~wire_out_quotient[9] ,  divisor[8] ,  wire_7_7_8_8_remainter ,  wire_8_8_9_9_remainter ,  wire_8_07_08_curry ,  wire_8_08_09_curry );
	div_cell cas_8_7 ( ~wire_out_quotient[9] ,  divisor[7] ,  wire_7_6_8_7_remainter ,  wire_8_7_9_8_remainter ,  wire_8_06_07_curry ,  wire_8_07_08_curry );
	div_cell cas_8_6 ( ~wire_out_quotient[9] ,  divisor[6] ,  wire_7_5_8_6_remainter ,  wire_8_6_9_7_remainter ,  wire_8_05_06_curry ,  wire_8_06_07_curry );
	div_cell cas_8_5 ( ~wire_out_quotient[9] ,  divisor[5] ,  wire_7_4_8_5_remainter ,  wire_8_5_9_6_remainter ,  wire_8_04_05_curry ,  wire_8_05_06_curry );
	div_cell cas_8_4 ( ~wire_out_quotient[9] ,  divisor[4] ,  wire_7_3_8_4_remainter ,  wire_8_4_9_5_remainter ,  wire_8_03_04_curry ,  wire_8_04_05_curry );
	div_cell cas_8_3 ( ~wire_out_quotient[9] ,  divisor[3] ,  wire_7_2_8_3_remainter ,  wire_8_3_9_4_remainter ,  wire_8_02_03_curry ,  wire_8_03_04_curry );
	div_cell cas_8_2 ( ~wire_out_quotient[9] ,  divisor[2] ,  wire_7_1_8_2_remainter ,  wire_8_2_9_3_remainter ,  wire_8_01_02_curry ,  wire_8_02_03_curry );
	div_cell cas_8_1 ( ~wire_out_quotient[9] ,  divisor[1] ,  wire_7_0_8_1_remainter ,  wire_8_1_9_2_remainter ,  wire_8_00_01_curry ,  wire_8_01_02_curry );
	
	div_cell cas_8_0 ( ~wire_out_quotient[9] ,  divisor[0] ,  dividend[8] ,  wire_8_0_9_1_remainter ,  ~wire_out_quotient[9] ,  wire_8_00_01_curry );

	//10th row
	div_cell cas_9_15 ( ~wire_out_quotient[8] ,  divisor[15] ,  wire_8_14_9_15_remainter ,   wire_out_quotient[7] ,  wire_9_14_15_curry ,  hang_9_wire_15 );

	div_cell cas_9_14 ( ~wire_out_quotient[8] ,  divisor[14] ,  wire_8_13_9_14_remainter ,  wire_9_14_10_15_remainter ,  wire_9_13_14_curry ,  wire_9_14_15_curry );
	div_cell cas_9_13 ( ~wire_out_quotient[8] ,  divisor[13] ,  wire_8_12_9_13_remainter ,  wire_9_13_10_14_remainter ,  wire_9_12_13_curry ,  wire_9_13_14_curry );
	div_cell cas_9_12 ( ~wire_out_quotient[8] ,  divisor[12] ,  wire_8_11_9_12_remainter ,  wire_9_12_10_13_remainter ,  wire_9_11_12_curry ,  wire_9_12_13_curry );
	div_cell cas_9_11 ( ~wire_out_quotient[8] ,  divisor[11] ,  wire_8_10_9_11_remainter ,  wire_9_11_10_12_remainter ,  wire_9_10_11_curry ,  wire_9_11_12_curry );
	div_cell cas_9_10 ( ~wire_out_quotient[8] ,  divisor[10] ,  wire_8_9_9_10_remainter ,  wire_9_10_10_11_remainter ,  wire_9_09_10_curry ,  wire_9_10_11_curry );
	div_cell cas_9_9 ( ~wire_out_quotient[8] ,  divisor[9] ,  wire_8_8_9_9_remainter ,  wire_9_9_10_10_remainter ,  wire_9_08_09_curry ,  wire_9_09_10_curry );
	div_cell cas_9_8 ( ~wire_out_quotient[8] ,  divisor[8] ,  wire_8_7_9_8_remainter ,  wire_9_8_10_9_remainter ,  wire_9_07_08_curry ,  wire_9_08_09_curry );
	div_cell cas_9_7 ( ~wire_out_quotient[8] ,  divisor[7] ,  wire_8_6_9_7_remainter ,  wire_9_7_10_8_remainter ,  wire_9_06_07_curry ,  wire_9_07_08_curry );
	div_cell cas_9_6 ( ~wire_out_quotient[8] ,  divisor[6] ,  wire_8_5_9_6_remainter ,  wire_9_6_10_7_remainter ,  wire_9_05_06_curry ,  wire_9_06_07_curry );
	div_cell cas_9_5 ( ~wire_out_quotient[8] ,  divisor[5] ,  wire_8_4_9_5_remainter ,  wire_9_5_10_6_remainter ,  wire_9_04_05_curry ,  wire_9_05_06_curry );
	div_cell cas_9_4 ( ~wire_out_quotient[8] ,  divisor[4] ,  wire_8_3_9_4_remainter ,  wire_9_4_10_5_remainter ,  wire_9_03_04_curry ,  wire_9_04_05_curry );
	div_cell cas_9_3 ( ~wire_out_quotient[8] ,  divisor[3] ,  wire_8_2_9_3_remainter ,  wire_9_3_10_4_remainter ,  wire_9_02_03_curry ,  wire_9_03_04_curry );
	div_cell cas_9_2 ( ~wire_out_quotient[8] ,  divisor[2] ,  wire_8_1_9_2_remainter ,  wire_9_2_10_3_remainter ,  wire_9_01_02_curry ,  wire_9_02_03_curry );
	div_cell cas_9_1 ( ~wire_out_quotient[8] ,  divisor[1] ,  wire_8_0_9_1_remainter ,  wire_9_1_10_2_remainter ,  wire_9_00_01_curry ,  wire_9_01_02_curry );
	
	div_cell cas_9_0 ( ~wire_out_quotient[8] ,  divisor[0] ,  dividend[7] ,  wire_9_0_10_1_remainter ,  ~wire_out_quotient[8] ,  wire_9_00_01_curry );

	//11th row
	div_cell cas_10_15 ( ~wire_out_quotient[7] ,  divisor[15] ,  wire_9_14_10_15_remainter ,   wire_out_quotient[6] ,  wire_10_14_15_curry ,  hang_10_wire_15 );

	div_cell cas_10_14 ( ~wire_out_quotient[7] ,  divisor[14] ,  wire_9_13_10_14_remainter ,  wire_10_14_11_15_remainter ,  wire_10_13_14_curry ,  wire_10_14_15_curry );
	div_cell cas_10_13 ( ~wire_out_quotient[7] ,  divisor[13] ,  wire_9_12_10_13_remainter ,  wire_10_13_11_14_remainter ,  wire_10_12_13_curry ,  wire_10_13_14_curry );
	div_cell cas_10_12 ( ~wire_out_quotient[7] ,  divisor[12] ,  wire_9_11_10_12_remainter ,  wire_10_12_11_13_remainter ,  wire_10_11_12_curry ,  wire_10_12_13_curry );
	div_cell cas_10_11 ( ~wire_out_quotient[7] ,  divisor[11] ,  wire_9_10_10_11_remainter ,  wire_10_11_11_12_remainter ,  wire_10_10_11_curry ,  wire_10_11_12_curry );
	div_cell cas_10_10 ( ~wire_out_quotient[7] ,  divisor[10] ,  wire_9_9_10_10_remainter ,  wire_10_10_11_11_remainter ,  wire_10_09_10_curry ,  wire_10_10_11_curry );
	div_cell cas_10_9 ( ~wire_out_quotient[7] ,  divisor[9] ,  wire_9_8_10_9_remainter ,  wire_10_9_11_10_remainter ,  wire_10_08_09_curry ,  wire_10_09_10_curry );
	div_cell cas_10_8 ( ~wire_out_quotient[7] ,  divisor[8] ,  wire_9_7_10_8_remainter ,  wire_10_8_11_9_remainter ,  wire_10_07_08_curry ,  wire_10_08_09_curry );
	div_cell cas_10_7 ( ~wire_out_quotient[7] ,  divisor[7] ,  wire_9_6_10_7_remainter ,  wire_10_7_11_8_remainter ,  wire_10_06_07_curry ,  wire_10_07_08_curry );
	div_cell cas_10_6 ( ~wire_out_quotient[7] ,  divisor[6] ,  wire_9_5_10_6_remainter ,  wire_10_6_11_7_remainter ,  wire_10_05_06_curry ,  wire_10_06_07_curry );
	div_cell cas_10_5 ( ~wire_out_quotient[7] ,  divisor[5] ,  wire_9_4_10_5_remainter ,  wire_10_5_11_6_remainter ,  wire_10_04_05_curry ,  wire_10_05_06_curry );
	div_cell cas_10_4 ( ~wire_out_quotient[7] ,  divisor[4] ,  wire_9_3_10_4_remainter ,  wire_10_4_11_5_remainter ,  wire_10_03_04_curry ,  wire_10_04_05_curry );
	div_cell cas_10_3 ( ~wire_out_quotient[7] ,  divisor[3] ,  wire_9_2_10_3_remainter ,  wire_10_3_11_4_remainter ,  wire_10_02_03_curry ,  wire_10_03_04_curry );
	div_cell cas_10_2 ( ~wire_out_quotient[7] ,  divisor[2] ,  wire_9_1_10_2_remainter ,  wire_10_2_11_3_remainter ,  wire_10_01_02_curry ,  wire_10_02_03_curry );
	div_cell cas_10_1 ( ~wire_out_quotient[7] ,  divisor[1] ,  wire_9_0_10_1_remainter ,  wire_10_1_11_2_remainter ,  wire_10_00_01_curry ,  wire_10_01_02_curry );
	
	div_cell cas_10_0 ( ~wire_out_quotient[7] ,  divisor[0] ,  dividend[6] ,  wire_10_0_11_1_remainter ,  ~wire_out_quotient[7] ,  wire_10_00_01_curry );

	//12th row
	div_cell cas_11_15 ( ~wire_out_quotient[6] ,  divisor[15] ,  wire_10_14_11_15_remainter ,   wire_out_quotient[5] ,  wire_11_14_15_curry ,  hang_11_wire_15 );

	div_cell cas_11_14 ( ~wire_out_quotient[6] ,  divisor[14] ,  wire_10_13_11_14_remainter ,  wire_11_14_12_15_remainter ,  wire_11_13_14_curry ,  wire_11_14_15_curry );
	div_cell cas_11_13 ( ~wire_out_quotient[6] ,  divisor[13] ,  wire_10_12_11_13_remainter ,  wire_11_13_12_14_remainter ,  wire_11_12_13_curry ,  wire_11_13_14_curry );
	div_cell cas_11_12 ( ~wire_out_quotient[6] ,  divisor[12] ,  wire_10_11_11_12_remainter ,  wire_11_12_12_13_remainter ,  wire_11_11_12_curry ,  wire_11_12_13_curry );
	div_cell cas_11_11 ( ~wire_out_quotient[6] ,  divisor[11] ,  wire_10_10_11_11_remainter ,  wire_11_11_12_12_remainter ,  wire_11_10_11_curry ,  wire_11_11_12_curry );
	div_cell cas_11_10 ( ~wire_out_quotient[6] ,  divisor[10] ,  wire_10_9_11_10_remainter ,  wire_11_10_12_11_remainter ,  wire_11_09_10_curry ,  wire_11_10_11_curry );
	div_cell cas_11_9 ( ~wire_out_quotient[6] ,  divisor[9] ,  wire_10_8_11_9_remainter ,  wire_11_9_12_10_remainter ,  wire_11_08_09_curry ,  wire_11_09_10_curry );
	div_cell cas_11_8 ( ~wire_out_quotient[6] ,  divisor[8] ,  wire_10_7_11_8_remainter ,  wire_11_8_12_9_remainter ,  wire_11_07_08_curry ,  wire_11_08_09_curry );
	div_cell cas_11_7 ( ~wire_out_quotient[6] ,  divisor[7] ,  wire_10_6_11_7_remainter ,  wire_11_7_12_8_remainter ,  wire_11_06_07_curry ,  wire_11_07_08_curry );
	div_cell cas_11_6 ( ~wire_out_quotient[6] ,  divisor[6] ,  wire_10_5_11_6_remainter ,  wire_11_6_12_7_remainter ,  wire_11_05_06_curry ,  wire_11_06_07_curry );
	div_cell cas_11_5 ( ~wire_out_quotient[6] ,  divisor[5] ,  wire_10_4_11_5_remainter ,  wire_11_5_12_6_remainter ,  wire_11_04_05_curry ,  wire_11_05_06_curry );
	div_cell cas_11_4 ( ~wire_out_quotient[6] ,  divisor[4] ,  wire_10_3_11_4_remainter ,  wire_11_4_12_5_remainter ,  wire_11_03_04_curry ,  wire_11_04_05_curry );
	div_cell cas_11_3 ( ~wire_out_quotient[6] ,  divisor[3] ,  wire_10_2_11_3_remainter ,  wire_11_3_12_4_remainter ,  wire_11_02_03_curry ,  wire_11_03_04_curry );
	div_cell cas_11_2 ( ~wire_out_quotient[6] ,  divisor[2] ,  wire_10_1_11_2_remainter ,  wire_11_2_12_3_remainter ,  wire_11_01_02_curry ,  wire_11_02_03_curry );
	div_cell cas_11_1 ( ~wire_out_quotient[6] ,  divisor[1] ,  wire_10_0_11_1_remainter ,  wire_11_1_12_2_remainter ,  wire_11_00_01_curry ,  wire_11_01_02_curry );
	
	div_cell cas_11_0 ( ~wire_out_quotient[6] ,  divisor[0] ,  dividend[5] ,  wire_11_0_12_1_remainter ,  ~wire_out_quotient[6] ,  wire_11_00_01_curry );

	//13th row
	div_cell cas_12_15 ( ~wire_out_quotient[5] ,  divisor[15] ,  wire_11_14_12_15_remainter ,   wire_out_quotient[4] ,  wire_12_14_15_curry ,  hang_12_wire_15 );
	div_cell cas_12_14 ( ~wire_out_quotient[5] ,  divisor[14] ,  wire_11_13_12_14_remainter ,  wire_12_14_13_15_remainter ,  wire_12_13_14_curry ,  wire_12_14_15_curry );
	div_cell cas_12_13 ( ~wire_out_quotient[5] ,  divisor[13] ,  wire_11_12_12_13_remainter ,  wire_12_13_13_14_remainter ,  wire_12_12_13_curry ,  wire_12_13_14_curry );
	div_cell cas_12_12 ( ~wire_out_quotient[5] ,  divisor[12] ,  wire_11_11_12_12_remainter ,  wire_12_12_13_13_remainter ,  wire_12_11_12_curry ,  wire_12_12_13_curry );
	div_cell cas_12_11 ( ~wire_out_quotient[5] ,  divisor[11] ,  wire_11_10_12_11_remainter ,  wire_12_11_13_12_remainter ,  wire_12_10_11_curry ,  wire_12_11_12_curry );
	div_cell cas_12_10 ( ~wire_out_quotient[5] ,  divisor[10] ,  wire_11_9_12_10_remainter ,  wire_12_10_13_11_remainter ,  wire_12_09_10_curry ,  wire_12_10_11_curry );
	div_cell cas_12_9 ( ~wire_out_quotient[5] ,  divisor[9] ,  wire_11_8_12_9_remainter ,  wire_12_9_13_10_remainter ,  wire_12_08_09_curry ,  wire_12_09_10_curry );
	div_cell cas_12_8 ( ~wire_out_quotient[5] ,  divisor[8] ,  wire_11_7_12_8_remainter ,  wire_12_8_13_9_remainter ,  wire_12_07_08_curry ,  wire_12_08_09_curry );
	div_cell cas_12_7 ( ~wire_out_quotient[5] ,  divisor[7] ,  wire_11_6_12_7_remainter ,  wire_12_7_13_8_remainter ,  wire_12_06_07_curry ,  wire_12_07_08_curry );
	div_cell cas_12_6 ( ~wire_out_quotient[5] ,  divisor[6] ,  wire_11_5_12_6_remainter ,  wire_12_6_13_7_remainter ,  wire_12_05_06_curry ,  wire_12_06_07_curry );
	div_cell cas_12_5 ( ~wire_out_quotient[5] ,  divisor[5] ,  wire_11_4_12_5_remainter ,  wire_12_5_13_6_remainter ,  wire_12_04_05_curry ,  wire_12_05_06_curry );
	div_cell cas_12_4 ( ~wire_out_quotient[5] ,  divisor[4] ,  wire_11_3_12_4_remainter ,  wire_12_4_13_5_remainter ,  wire_12_03_04_curry ,  wire_12_04_05_curry );
	div_cell cas_12_3 ( ~wire_out_quotient[5] ,  divisor[3] ,  wire_11_2_12_3_remainter ,  wire_12_3_13_4_remainter ,  wire_12_02_03_curry ,  wire_12_03_04_curry );
	div_cell cas_12_2 ( ~wire_out_quotient[5] ,  divisor[2] ,  wire_11_1_12_2_remainter ,  wire_12_2_13_3_remainter ,  wire_12_01_02_curry ,  wire_12_02_03_curry );
	div_cell cas_12_1 ( ~wire_out_quotient[5] ,  divisor[1] ,  wire_11_0_12_1_remainter ,  wire_12_1_13_2_remainter ,  wire_12_00_01_curry ,  wire_12_01_02_curry );
	
	div_cell cas_12_0 ( ~wire_out_quotient[5] ,  divisor[0] ,  dividend[4] ,  wire_12_0_13_1_remainter ,  ~wire_out_quotient[5] ,  wire_12_00_01_curry );

	//14th row
	div_cell cas_13_15 ( ~wire_out_quotient[4] ,  divisor[15] ,  wire_12_14_13_15_remainter ,   wire_out_quotient[3] ,  wire_13_14_15_curry ,  hang_13_wire_15 );

	div_cell cas_13_14 ( ~wire_out_quotient[4] ,  divisor[14] ,  wire_12_13_13_14_remainter ,  wire_13_14_14_15_remainter ,  wire_13_13_14_curry ,  wire_13_14_15_curry );
	div_cell cas_13_13 ( ~wire_out_quotient[4] ,  divisor[13] ,  wire_12_12_13_13_remainter ,  wire_13_13_14_14_remainter ,  wire_13_12_13_curry ,  wire_13_13_14_curry );
	div_cell cas_13_12 ( ~wire_out_quotient[4] ,  divisor[12] ,  wire_12_11_13_12_remainter ,  wire_13_12_14_13_remainter ,  wire_13_11_12_curry ,  wire_13_12_13_curry );
	div_cell cas_13_11 ( ~wire_out_quotient[4] ,  divisor[11] ,  wire_12_10_13_11_remainter ,  wire_13_11_14_12_remainter ,  wire_13_10_11_curry ,  wire_13_11_12_curry );
	div_cell cas_13_10 ( ~wire_out_quotient[4] ,  divisor[10] ,  wire_12_9_13_10_remainter ,  wire_13_10_14_11_remainter ,  wire_13_09_10_curry ,  wire_13_10_11_curry );
	div_cell cas_13_9 ( ~wire_out_quotient[4] ,  divisor[9] ,  wire_12_8_13_9_remainter ,  wire_13_9_14_10_remainter ,  wire_13_08_09_curry ,  wire_13_09_10_curry );
	div_cell cas_13_8 ( ~wire_out_quotient[4] ,  divisor[8] ,  wire_12_7_13_8_remainter ,  wire_13_8_14_9_remainter ,  wire_13_07_08_curry ,  wire_13_08_09_curry );
	div_cell cas_13_7 ( ~wire_out_quotient[4] ,  divisor[7] ,  wire_12_6_13_7_remainter ,  wire_13_7_14_8_remainter ,  wire_13_06_07_curry ,  wire_13_07_08_curry );
	div_cell cas_13_6 ( ~wire_out_quotient[4] ,  divisor[6] ,  wire_12_5_13_6_remainter ,  wire_13_6_14_7_remainter ,  wire_13_05_06_curry ,  wire_13_06_07_curry );
	div_cell cas_13_5 ( ~wire_out_quotient[4] ,  divisor[5] ,  wire_12_4_13_5_remainter ,  wire_13_5_14_6_remainter ,  wire_13_04_05_curry ,  wire_13_05_06_curry );
	div_cell cas_13_4 ( ~wire_out_quotient[4] ,  divisor[4] ,  wire_12_3_13_4_remainter ,  wire_13_4_14_5_remainter ,  wire_13_03_04_curry ,  wire_13_04_05_curry );
	div_cell cas_13_3 ( ~wire_out_quotient[4] ,  divisor[3] ,  wire_12_2_13_3_remainter ,  wire_13_3_14_4_remainter ,  wire_13_02_03_curry ,  wire_13_03_04_curry );
	div_cell cas_13_2 ( ~wire_out_quotient[4] ,  divisor[2] ,  wire_12_1_13_2_remainter ,  wire_13_2_14_3_remainter ,  wire_13_01_02_curry ,  wire_13_02_03_curry );
	div_cell cas_13_1 ( ~wire_out_quotient[4] ,  divisor[1] ,  wire_12_0_13_1_remainter ,  wire_13_1_14_2_remainter ,  wire_13_00_01_curry ,  wire_13_01_02_curry );
	
	div_cell cas_13_0 ( ~wire_out_quotient[4] ,  divisor[0] ,  dividend[3] ,  wire_13_0_14_1_remainter ,  ~wire_out_quotient[4] ,  wire_13_00_01_curry );

	//15th row
	div_cell cas_14_15 ( ~wire_out_quotient[3] ,  divisor[15] ,  wire_13_14_14_15_remainter ,   wire_out_quotient[2] ,  wire_14_14_15_curry ,  hang_14_wire_15 );

	div_cell cas_14_14 ( ~wire_out_quotient[3] ,  divisor[14] ,  wire_13_13_14_14_remainter ,  wire_14_14_15_15_remainter ,  wire_14_13_14_curry ,  wire_14_14_15_curry );
	div_cell cas_14_13 ( ~wire_out_quotient[3] ,  divisor[13] ,  wire_13_12_14_13_remainter ,  wire_14_13_15_14_remainter ,  wire_14_12_13_curry ,  wire_14_13_14_curry );
	div_cell cas_14_12 ( ~wire_out_quotient[3] ,  divisor[12] ,  wire_13_11_14_12_remainter ,  wire_14_12_15_13_remainter ,  wire_14_11_12_curry ,  wire_14_12_13_curry );
	div_cell cas_14_11 ( ~wire_out_quotient[3] ,  divisor[11] ,  wire_13_10_14_11_remainter ,  wire_14_11_15_12_remainter ,  wire_14_10_11_curry ,  wire_14_11_12_curry );
	div_cell cas_14_10 ( ~wire_out_quotient[3] ,  divisor[10] ,  wire_13_9_14_10_remainter ,  wire_14_10_15_11_remainter ,  wire_14_09_10_curry ,  wire_14_10_11_curry );
	div_cell cas_14_9 ( ~wire_out_quotient[3] ,  divisor[9] ,  wire_13_8_14_9_remainter ,  wire_14_9_15_10_remainter ,  wire_14_08_09_curry ,  wire_14_09_10_curry );
	div_cell cas_14_8 ( ~wire_out_quotient[3] ,  divisor[8] ,  wire_13_7_14_8_remainter ,  wire_14_8_15_9_remainter ,  wire_14_07_08_curry ,  wire_14_08_09_curry );
	div_cell cas_14_7 ( ~wire_out_quotient[3] ,  divisor[7] ,  wire_13_6_14_7_remainter ,  wire_14_7_15_8_remainter ,  wire_14_06_07_curry ,  wire_14_07_08_curry );
	div_cell cas_14_6 ( ~wire_out_quotient[3] ,  divisor[6] ,  wire_13_5_14_6_remainter ,  wire_14_6_15_7_remainter ,  wire_14_05_06_curry ,  wire_14_06_07_curry );
	div_cell cas_14_5 ( ~wire_out_quotient[3] ,  divisor[5] ,  wire_13_4_14_5_remainter ,  wire_14_5_15_6_remainter ,  wire_14_04_05_curry ,  wire_14_05_06_curry );
	div_cell cas_14_4 ( ~wire_out_quotient[3] ,  divisor[4] ,  wire_13_3_14_4_remainter ,  wire_14_4_15_5_remainter ,  wire_14_03_04_curry ,  wire_14_04_05_curry );
	div_cell cas_14_3 ( ~wire_out_quotient[3] ,  divisor[3] ,  wire_13_2_14_3_remainter ,  wire_14_3_15_4_remainter ,  wire_14_02_03_curry ,  wire_14_03_04_curry );
	div_cell cas_14_2 ( ~wire_out_quotient[3] ,  divisor[2] ,  wire_13_1_14_2_remainter ,  wire_14_2_15_3_remainter ,  wire_14_01_02_curry ,  wire_14_02_03_curry );
	div_cell cas_14_1 ( ~wire_out_quotient[3] ,  divisor[1] ,  wire_13_0_14_1_remainter ,  wire_14_1_15_2_remainter ,  wire_14_00_01_curry ,  wire_14_01_02_curry );
	
	div_cell cas_14_0 ( ~wire_out_quotient[3] ,  divisor[0] ,  dividend[2] ,  wire_14_0_15_1_remainter ,  ~wire_out_quotient[3] ,  wire_14_00_01_curry );

	//16th row
	div_cell cas_15_15 ( ~wire_out_quotient[2] ,  divisor[15] ,  wire_14_14_15_15_remainter ,   wire_out_quotient[1] ,  wire_15_14_15_curry ,  hang_15_wire_15 );

	div_cell cas_15_14 ( ~wire_out_quotient[2] ,  divisor[14] ,  wire_14_13_15_14_remainter ,  wire_15_14_16_15_remainter ,  wire_15_13_14_curry ,  wire_15_14_15_curry );
	div_cell cas_15_13 ( ~wire_out_quotient[2] ,  divisor[13] ,  wire_14_12_15_13_remainter ,  wire_15_13_16_14_remainter ,  wire_15_12_13_curry ,  wire_15_13_14_curry );
	div_cell cas_15_12 ( ~wire_out_quotient[2] ,  divisor[12] ,  wire_14_11_15_12_remainter ,  wire_15_12_16_13_remainter ,  wire_15_11_12_curry ,  wire_15_12_13_curry );
	div_cell cas_15_11 ( ~wire_out_quotient[2] ,  divisor[11] ,  wire_14_10_15_11_remainter ,  wire_15_11_16_12_remainter ,  wire_15_10_11_curry ,  wire_15_11_12_curry );
	div_cell cas_15_10 ( ~wire_out_quotient[2] ,  divisor[10] ,  wire_14_9_15_10_remainter ,  wire_15_10_16_11_remainter ,  wire_15_09_10_curry ,  wire_15_10_11_curry );
	div_cell cas_15_9 ( ~wire_out_quotient[2] ,  divisor[9] ,  wire_14_8_15_9_remainter ,  wire_15_9_16_10_remainter ,  wire_15_08_09_curry ,  wire_15_09_10_curry );
	div_cell cas_15_8 ( ~wire_out_quotient[2] ,  divisor[8] ,  wire_14_7_15_8_remainter ,  wire_15_8_16_9_remainter ,  wire_15_07_08_curry ,  wire_15_08_09_curry );
	div_cell cas_15_7 ( ~wire_out_quotient[2] ,  divisor[7] ,  wire_14_6_15_7_remainter ,  wire_15_7_16_8_remainter ,  wire_15_06_07_curry ,  wire_15_07_08_curry );
	div_cell cas_15_6 ( ~wire_out_quotient[2] ,  divisor[6] ,  wire_14_5_15_6_remainter ,  wire_15_6_16_7_remainter ,  wire_15_05_06_curry ,  wire_15_06_07_curry );
	div_cell cas_15_5 ( ~wire_out_quotient[2] ,  divisor[5] ,  wire_14_4_15_5_remainter ,  wire_15_5_16_6_remainter ,  wire_15_04_05_curry ,  wire_15_05_06_curry );
	div_cell cas_15_4 ( ~wire_out_quotient[2] ,  divisor[4] ,  wire_14_3_15_4_remainter ,  wire_15_4_16_5_remainter ,  wire_15_03_04_curry ,  wire_15_04_05_curry );
	div_cell cas_15_3 ( ~wire_out_quotient[2] ,  divisor[3] ,  wire_14_2_15_3_remainter ,  wire_15_3_16_4_remainter ,  wire_15_02_03_curry ,  wire_15_03_04_curry );
	div_cell cas_15_2 ( ~wire_out_quotient[2] ,  divisor[2] ,  wire_14_1_15_2_remainter ,  wire_15_2_16_3_remainter ,  wire_15_01_02_curry ,  wire_15_02_03_curry );
	div_cell cas_15_1 ( ~wire_out_quotient[2] ,  divisor[1] ,  wire_14_0_15_1_remainter ,  wire_15_1_16_2_remainter ,  wire_15_00_01_curry ,  wire_15_01_02_curry );
	
	div_cell cas_15_0 ( ~wire_out_quotient[2] ,  divisor[0] ,  dividend[1] ,  wire_15_0_16_1_remainter ,  ~wire_out_quotient[2] ,  wire_15_00_01_curry );

	//17th row
	div_cell cas_16_15 ( ~wire_out_quotient[1] ,  divisor[15] ,  wire_15_14_16_15_remainter ,   wire_out_quotient[0] ,  wire_16_14_15_curry ,  hang_16_wire_15 );

	div_cell cas_16_14 ( ~wire_out_quotient[1] ,  divisor[14] ,  wire_15_13_16_14_remainter ,  wire_out_remainder[14] ,  wire_16_13_14_curry ,  wire_16_14_15_curry );
	div_cell cas_16_13 ( ~wire_out_quotient[1] ,  divisor[13] ,  wire_15_12_16_13_remainter ,  wire_out_remainder[13] ,  wire_16_12_13_curry ,  wire_16_13_14_curry );
	div_cell cas_16_12 ( ~wire_out_quotient[1] ,  divisor[12] ,  wire_15_11_16_12_remainter ,  wire_out_remainder[12] ,  wire_16_11_12_curry ,  wire_16_12_13_curry );
	div_cell cas_16_11 ( ~wire_out_quotient[1] ,  divisor[11] ,  wire_15_10_16_11_remainter ,  wire_out_remainder[11] ,  wire_16_10_11_curry ,  wire_16_11_12_curry );
	div_cell cas_16_10 ( ~wire_out_quotient[1] ,  divisor[10] ,  wire_15_9_16_10_remainter ,  wire_out_remainder[10] ,  wire_16_09_10_curry ,  wire_16_10_11_curry );
	div_cell cas_16_9 ( ~wire_out_quotient[1] ,  divisor[9] ,  wire_15_8_16_9_remainter ,  wire_out_remainder[9] ,  wire_16_08_09_curry ,  wire_16_09_10_curry );
	div_cell cas_16_8 ( ~wire_out_quotient[1] ,  divisor[8] ,  wire_15_7_16_8_remainter ,  wire_out_remainder[8] ,  wire_16_07_08_curry ,  wire_16_08_09_curry );
	div_cell cas_16_7 ( ~wire_out_quotient[1] ,  divisor[7] ,  wire_15_6_16_7_remainter ,  wire_out_remainder[7] ,  wire_16_06_07_curry ,  wire_16_07_08_curry );
	div_cell cas_16_6 ( ~wire_out_quotient[1] ,  divisor[6] ,  wire_15_5_16_6_remainter ,  wire_out_remainder[6] ,  wire_16_05_06_curry ,  wire_16_06_07_curry );
	div_cell cas_16_5 ( ~wire_out_quotient[1] ,  divisor[5] ,  wire_15_4_16_5_remainter ,  wire_out_remainder[5] ,  wire_16_04_05_curry ,  wire_16_05_06_curry );
	div_cell cas_16_4 ( ~wire_out_quotient[1] ,  divisor[4] ,  wire_15_3_16_4_remainter ,  wire_out_remainder[4] ,  wire_16_03_04_curry ,  wire_16_04_05_curry );
	div_cell cas_16_3 ( ~wire_out_quotient[1] ,  divisor[3] ,  wire_15_2_16_3_remainter ,  wire_out_remainder[3] ,  wire_16_02_03_curry ,  wire_16_03_04_curry );
	div_cell cas_16_2 ( ~wire_out_quotient[1] ,  divisor[2] ,  wire_15_1_16_2_remainter ,  wire_out_remainder[2] ,  wire_16_01_02_curry ,  wire_16_02_03_curry );
	div_cell cas_16_1 ( ~wire_out_quotient[1] ,  divisor[1] ,  wire_15_0_16_1_remainter ,  wire_out_remainder[1] ,  wire_16_00_01_curry ,  wire_16_01_02_curry );
	
	div_cell cas_16_0 ( ~wire_out_quotient[1] ,  divisor[0] ,  dividend[0] ,  wire_out_remainder[0] ,  ~wire_out_quotient[1] ,  wire_16_00_01_curry );

endmodule // interconect_cells