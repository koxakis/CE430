module interconect_cells(
	clk,
	reset,
	divisor,
	dividend,
	mode,
	valid_input,
	valid_output,
	final_output
);

	input [31:0] dividend;
	input [15:0] divisor;

	input clk, reset;
	input valid_input;

	output valid_output;
	output [16:0] final_output;

	assign final_output = (mode) div_res : mod_res;

	assign div_res[15] = ~wire_out_quotient_15;
	assign div_res[14] = ~wire_out_quotient_14;
	assign div_res[13] = ~wire_out_quotient_13;
	assign div_res[12] = ~wire_out_quotient_12;
	assign div_res[11] = ~wire_out_quotient_11;
	assign div_res[10] = ~wire_out_quotient_10;
	assign div_res[9] = ~wire_out_quotient_9;
	assign div_res[8] = ~wire_out_quotient_8;
	assign div_res[7] = ~wire_out_quotient_7;
	assign div_res[6] = ~wire_out_quotient_6;
	assign div_res[5] = ~wire_out_quotient_5;
	assign div_res[4] = ~wire_out_quotient_4;
	assign div_res[3] = ~wire_out_quotient_3;
	assign div_res[2] = ~wire_out_quotient_2;
	assign div_res[1] = ~wire_out_quotient_1;
	assign div_res[0] = ~wire_out_quotient_0;

	assign mod_res[14] = wire_out_remainder_15;
	assign mod_res[14] = wire_out_remainder_14;
	assign mod_res[13] = wire_out_remainder_13;
	assign mod_res[12] = wire_out_remainder_12;
	assign mod_res[11] = wire_out_remainder_11;
	assign mod_res[10] = wire_out_remainder_10;
	assign mod_res[9] = wire_out_remainder_9;
	assign mod_res[8] = wire_out_remainder_8;
	assign mod_res[7] = wire_out_remainder_7;
	assign mod_res[6] = wire_out_remainder_6;
	assign mod_res[5] = wire_out_remainder_5;
	assign mod_res[4] = wire_out_remainder_4;
	assign mod_res[3] = wire_out_remainder_3;
	assign mod_res[2] = wire_out_remainder_2;
	assign mod_res[1] = wire_out_remainder_1;
	assign mod_res[0] = wire_out_remainder_0;	

	//div_cell cas_X_Y (T_in,Divisor_in,Remainder_in/dividend,Remainder_out,C_in,C_out);
	//. (T_in), . (Divisor_in), . (Remainder_in), . (Remainder_out), . (C_in), . (C_out)
	//1st row
	div_cell cas_0_15 (.1'b1(T_in), .divisor[15](Divisor_in), .dividend[31](Remainder_in), .wire_out_quotient_15(Remainder_out), .wire_0_14_15_curry(C_in), .hang_0_wire_15(C_out));

	div_cell cas_0_14 (.1'b1(T_in), .divisor[14](Divisor_in), .dividend[30](Remainder_in), .wire_0_14_1_15_remainter(Remainder_out), .wire_0_13_14_curry(C_in), .wire_0_14_15_curry(C_out));
	div_cell cas_0_13 (.1'b1(T_in), .divisor[13](Divisor_in), .dividend[29](Remainder_in), .wire_0_13_1_14_remainter(Remainder_out), .wire_0_12_13_curry(C_in), .wire_0_13_14_curry(C_out));
	div_cell cas_0_12 (.1'b1(T_in), .divisor[12](Divisor_in), .dividend[28](Remainder_in), .wire_0_12_1_13_remainter(Remainder_out), .wire_0_11_12_curry(C_in), .wire_0_12_13_curry(C_out));
	div_cell cas_0_11 (.1'b1(T_in), .divisor[11](Divisor_in), .dividend[27](Remainder_in), .wire_0_11_1_12_remainter(Remainder_out), .wire_0_10_11_curry(C_in), .wire_0_11_12_curry(C_out));
	div_cell cas_0_10 (.1'b1(T_in), .divisor[10](Divisor_in), .dividend[26](Remainder_in), .wire_0_10_1_11_remainter(Remainder_out), .wire_0_09_10_curry(C_in), .wire_0_10_11_curry(C_out));
	div_cell cas_0_9 (.1'b1(T_in), .divisor[9](Divisor_in), .dividend[25](Remainder_in), .wire_0_9_1_10_remainter(Remainder_out), .wire_0_08_09_curry(C_in), .wire_0_09_10_curry(C_out));
	div_cell cas_0_8 (.1'b1(T_in), .divisor[8](Divisor_in), .dividend[24](Remainder_in), .wire_0_8_1_9_remainter(Remainder_out), .wire_0_07_08_curry(C_in), .wire_0_08_09_curry(C_out));
	div_cell cas_0_7 (.1'b1(T_in), .divisor[7](Divisor_in), .dividend[23](Remainder_in), .wire_0_7_1_8_remainter(Remainder_out), .wire_0_06_07_curry(C_in), .wire_0_07_08_curry(C_out));
	div_cell cas_0_6 (.1'b1(T_in), .divisor[6](Divisor_in), .dividend[22](Remainder_in), .wire_0_6_1_7_remainter(Remainder_out), .wire_0_05_06_curry(C_in), .wire_0_06_07_curry(C_out));
	div_cell cas_0_5 (.1'b1(T_in), .divisor[5](Divisor_in), .dividend[21](Remainder_in), .wire_0_5_1_6_remainter(Remainder_out), .wire_0_04_05_curry(C_in), .wire_0_05_06_curry(C_out));
	div_cell cas_0_4 (.1'b1(T_in), .divisor[4](Divisor_in), .dividend[20](Remainder_in), .wire_0_4_1_5_remainter(Remainder_out), .wire_0_03_04_curry(C_in), .wire_0_04_05_curry(C_out));
	div_cell cas_0_3 (.1'b1(T_in), .divisor[3](Divisor_in), .dividend[19](Remainder_in), .wire_0_3_1_4_remainter(Remainder_out), .wire_0_02_03_curry(C_in), .wire_0_03_04_curry(C_out));
	div_cell cas_0_2 (.1'b1(T_in), .divisor[2](Divisor_in), .dividend[18](Remainder_in), .wire_0_2_1_3_remainter(Remainder_out), .wire_0_01_02_curry(C_in), .wire_0_02_03_curry(C_out));
	div_cell cas_0_1 (.1'b1(T_in), .divisor[1](Divisor_in), .dividend[17](Remainder_in), .wire_0_1_1_2_remainter(Remainder_out), .wire_0_00_01_curry(C_in), .wire_0_01_02_curry(C_out));

	div_cell cas_0_0 (.1'b1(T_in), .divisor[0](Divisor_in), .dividend[16](Remainder_in), .wire_0_0_1_1_remainter(Remainder_out), .1'b1(C_in), .wire_0_00_01_curry(C_out));

	//div_cell cas_X_Y (T_in,Divisor_in,Remainder_in/dividend,Remainder_out,C_in,C_out);
	//. (T_in), . (Divisor_in), . (Remainder_in), . (Remainder_out), . (C_in), . (C_out)
	//2nd row
	div_cell cas_1_15 (.~wire_out_quotient_15(T_in), .divisor[15](Divisor_in), .wire_0_14_1_15_remainter(Remainder_in), .wire_out_quotient_14(Remainder_out), .wire_1_14_15_curry(C_in), .hang_1_wire_15(C_out));

	div_cell cas_1_14 (.~wire_out_quotient_15(T_in), .divisor[14](Divisor_in), .wire_0_13_1_14_remainter(Remainder_in), .wire_1_14_2_15_remainter(Remainder_out), .wire_1_13_14_curry(C_in), .wire_1_14_15_curry(C_out));
	div_cell cas_1_13 (.~wire_out_quotient_15(T_in), .divisor[13](Divisor_in), .wire_0_12_1_13_remainter(Remainder_in), .wire_1_13_2_14_remainter(Remainder_out), .wire_1_12_13_curry(C_in), .wire_1_13_14_curry(C_out));
	div_cell cas_1_12 (.~wire_out_quotient_15(T_in), .divisor[12](Divisor_in), .wire_0_11_1_12_remainter(Remainder_in), .wire_1_12_2_13_remainter(Remainder_out), .wire_1_11_12_curry(C_in), .wire_1_12_13_curry(C_out));
	div_cell cas_1_11 (.~wire_out_quotient_15(T_in), .divisor[11](Divisor_in), .wire_0_10_1_11_remainter(Remainder_in), .wire_1_11_2_12_remainter(Remainder_out), .wire_1_10_11_curry(C_in), .wire_1_11_12_curry(C_out));
	div_cell cas_1_10 (.~wire_out_quotient_15(T_in), .divisor[10](Divisor_in), .wire_0_9_1_10_remainter(Remainder_in), .wire_1_10_2_11_remainter(Remainder_out), .wire_1_09_10_curry(C_in), .wire_1_10_11_curry(C_out));
	div_cell cas_1_9 (.~wire_out_quotient_15(T_in), .divisor[9](Divisor_in), .wire_0_8_1_9_remainter(Remainder_in), .wire_1_9_2_10_remainter(Remainder_out), .wire_1_08_09_curry(C_in), .wire_1_09_10_curry(C_out));
	div_cell cas_1_8 (.~wire_out_quotient_15(T_in), .divisor[8](Divisor_in), .wire_0_7_1_8_remainter(Remainder_in), .wire_1_8_2_9_remainter(Remainder_out), .wire_1_07_08_curry(C_in), .wire_1_08_09_curry(C_out));
	div_cell cas_1_7 (.~wire_out_quotient_15(T_in), .divisor[7](Divisor_in), .wire_0_6_1_7_remainter(Remainder_in), .wire_1_7_2_8_remainter(Remainder_out), .wire_1_06_07_curry(C_in), .wire_1_07_08_curry(C_out));
	div_cell cas_1_6 (.~wire_out_quotient_15(T_in), .divisor[6](Divisor_in), .wire_0_5_1_6_remainter(Remainder_in), .wire_1_6_2_7_remainter(Remainder_out), .wire_1_05_06_curry(C_in), .wire_1_06_07_curry(C_out));
	div_cell cas_1_5 (.~wire_out_quotient_15(T_in), .divisor[5](Divisor_in), .wire_0_4_1_5_remainter(Remainder_in), .wire_1_5_2_6_remainter(Remainder_out), .wire_1_04_05_curry(C_in), .wire_1_05_06_curry(C_out));
	div_cell cas_1_4 (.~wire_out_quotient_15(T_in), .divisor[4](Divisor_in), .wire_0_3_1_4_remainter(Remainder_in), .wire_1_4_2_5_remainter(Remainder_out), .wire_1_03_04_curry(C_in), .wire_1_04_05_curry(C_out));
	div_cell cas_1_3 (.~wire_out_quotient_15(T_in), .divisor[3](Divisor_in), .wire_0_2_1_3_remainter(Remainder_in), .wire_1_3_2_4_remainter(Remainder_out), .wire_1_02_03_curry(C_in), .wire_1_03_04_curry(C_out));
	div_cell cas_1_2 (.~wire_out_quotient_15(T_in), .divisor[2](Divisor_in), .wire_0_1_1_2_remainter(Remainder_in), .wire_1_2_2_3_remainter(Remainder_out), .wire_1_01_02_curry(C_in), .wire_1_02_03_curry(C_out));
	div_cell cas_1_1 (.~wire_out_quotient_15(T_in), .divisor[1](Divisor_in), .wire_0_0_1_1_remainter(Remainder_in), .wire_1_1_2_2_remainter(Remainder_out), .wire_1_00_01_curry(C_in), .wire_1_01_02_curry(C_out));

	div_cell cas_1_0 (.~wire_out_quotient_15(T_in), .divisor[0](Divisor_in), .dividend[15](Remainder_in), .wire_1_0_2_1_remainter(Remainder_out), .~wire_out_quotient_15(C_in), .wire_1_00_01_curry(C_out));

	//3rd row
	div_cell cas_2_15 (.~wire_out_quotient_14(T_in), .divisor[15](Divisor_in), .wire_1_14_2_15_remainter(Remainder_in), .wire_out_quotient_13(Remainder_out), .wire_2_14_15_curry(C_in), .hang_2_wire_15(C_out));

	div_cell cas_2_14 (.~wire_out_quotient_14(T_in), .divisor[14](Divisor_in), .wire_1_13_2_14_remainter(Remainder_in), .wire_2_14_3_15_remainter(Remainder_out), .wire_2_13_14_curry(C_in), .wire_2_14_15_curry(C_out));
	div_cell cas_2_13 (.~wire_out_quotient_14(T_in), .divisor[13](Divisor_in), .wire_1_12_2_13_remainter(Remainder_in), .wire_2_13_3_14_remainter(Remainder_out), .wire_2_12_13_curry(C_in), .wire_2_13_14_curry(C_out));
	div_cell cas_2_12 (.~wire_out_quotient_14(T_in), .divisor[12](Divisor_in), .wire_1_11_2_12_remainter(Remainder_in), .wire_2_12_3_13_remainter(Remainder_out), .wire_2_11_12_curry(C_in), .wire_2_12_13_curry(C_out));
	div_cell cas_2_11 (.~wire_out_quotient_14(T_in), .divisor[11](Divisor_in), .wire_1_10_2_11_remainter(Remainder_in), .wire_2_11_3_12_remainter(Remainder_out), .wire_2_10_11_curry(C_in), .wire_2_11_12_curry(C_out));
	div_cell cas_2_10 (.~wire_out_quotient_14(T_in), .divisor[10](Divisor_in), .wire_1_9_2_10_remainter(Remainder_in), .wire_2_10_3_11_remainter(Remainder_out), .wire_2_09_10_curry(C_in), .wire_2_10_11_curry(C_out));
	div_cell cas_2_9 (.~wire_out_quotient_14(T_in), .divisor[9](Divisor_in), .wire_1_8_2_9_remainter(Remainder_in), .wire_2_9_3_10_remainter(Remainder_out), .wire_2_08_09_curry(C_in), .wire_2_09_10_curry(C_out));
	div_cell cas_2_8 (.~wire_out_quotient_14(T_in), .divisor[8](Divisor_in), .wire_1_7_2_8_remainter(Remainder_in), .wire_2_8_3_9_remainter(Remainder_out), .wire_2_07_08_curry(C_in), .wire_2_08_09_curry(C_out));
	div_cell cas_2_7 (.~wire_out_quotient_14(T_in), .divisor[7](Divisor_in), .wire_1_6_2_7_remainter(Remainder_in), .wire_2_7_3_8_remainter(Remainder_out), .wire_2_06_07_curry(C_in), .wire_2_07_08_curry(C_out));
	div_cell cas_2_6 (.~wire_out_quotient_14(T_in), .divisor[6](Divisor_in), .wire_1_5_2_6_remainter(Remainder_in), .wire_2_6_3_7_remainter(Remainder_out), .wire_2_05_06_curry(C_in), .wire_2_06_07_curry(C_out));
	div_cell cas_2_5 (.~wire_out_quotient_14(T_in), .divisor[5](Divisor_in), .wire_1_4_2_5_remainter(Remainder_in), .wire_2_5_3_6_remainter(Remainder_out), .wire_2_04_05_curry(C_in), .wire_2_05_06_curry(C_out));
	div_cell cas_2_4 (.~wire_out_quotient_14(T_in), .divisor[4](Divisor_in), .wire_1_3_2_4_remainter(Remainder_in), .wire_2_4_3_5_remainter(Remainder_out), .wire_2_03_04_curry(C_in), .wire_2_04_05_curry(C_out));
	div_cell cas_2_3 (.~wire_out_quotient_14(T_in), .divisor[3](Divisor_in), .wire_1_2_2_3_remainter(Remainder_in), .wire_2_3_3_4_remainter(Remainder_out), .wire_2_02_03_curry(C_in), .wire_2_03_04_curry(C_out));
	div_cell cas_2_2 (.~wire_out_quotient_14(T_in), .divisor[2](Divisor_in), .wire_1_1_2_2_remainter(Remainder_in), .wire_2_2_3_3_remainter(Remainder_out), .wire_2_01_02_curry(C_in), .wire_2_02_03_curry(C_out));
	div_cell cas_2_1 (.~wire_out_quotient_14(T_in), .divisor[1](Divisor_in), .wire_1_0_2_1_remainter(Remainder_in), .wire_2_1_3_2_remainter(Remainder_out), .wire_2_00_01_curry(C_in), .wire_2_01_02_curry(C_out));

	div_cell cas_2_0 (.~wire_out_quotient_14(T_in), .divisor[0](Divisor_in), .dividend[14](Remainder_in), .wire_2_0_3_1_remainter(Remainder_out), .~wire_out_quotient_14(C_in), .wire_2_00_01_curry(C_out));

	//4th row
	div_cell cas_3_15 (.~wire_out_quotient_13(T_in), .divisor[15](Divisor_in), .wire_2_14_3_15_remainter(Remainder_in), .wire_out_quotient_12(Remainder_out), .wire_3_14_15_curry(C_in), .hang_3_wire_15(C_out));

	div_cell cas_3_14 (.~wire_out_quotient_13(T_in), .divisor[14](Divisor_in), .wire_2_13_3_14_remainter(Remainder_in), .wire_3_14_4_15_remainter(Remainder_out), .wire_3_13_14_curry(C_in), .wire_3_14_15_curry(C_out));
	div_cell cas_3_13 (.~wire_out_quotient_13(T_in), .divisor[13](Divisor_in), .wire_2_12_3_13_remainter(Remainder_in), .wire_3_13_4_14_remainter(Remainder_out), .wire_3_12_13_curry(C_in), .wire_3_13_14_curry(C_out));
	div_cell cas_3_12 (.~wire_out_quotient_13(T_in), .divisor[12](Divisor_in), .wire_2_11_3_12_remainter(Remainder_in), .wire_3_12_4_13_remainter(Remainder_out), .wire_3_11_12_curry(C_in), .wire_3_12_13_curry(C_out));
	div_cell cas_3_11 (.~wire_out_quotient_13(T_in), .divisor[11](Divisor_in), .wire_2_10_3_11_remainter(Remainder_in), .wire_3_11_4_12_remainter(Remainder_out), .wire_3_10_11_curry(C_in), .wire_3_11_12_curry(C_out));
	div_cell cas_3_10 (.~wire_out_quotient_13(T_in), .divisor[10](Divisor_in), .wire_2_9_3_10_remainter(Remainder_in), .wire_3_10_4_11_remainter(Remainder_out), .wire_3_09_10_curry(C_in), .wire_3_10_11_curry(C_out));
	div_cell cas_3_9 (.~wire_out_quotient_13(T_in), .divisor[9](Divisor_in), .wire_2_8_3_9_remainter(Remainder_in), .wire_3_9_4_10_remainter(Remainder_out), .wire_3_08_09_curry(C_in), .wire_3_09_10_curry(C_out));
	div_cell cas_3_8 (.~wire_out_quotient_13(T_in), .divisor[8](Divisor_in), .wire_2_7_3_8_remainter(Remainder_in), .wire_3_8_4_9_remainter(Remainder_out), .wire_3_07_08_curry(C_in), .wire_3_08_09_curry(C_out));
	div_cell cas_3_7 (.~wire_out_quotient_13(T_in), .divisor[7](Divisor_in), .wire_2_6_3_7_remainter(Remainder_in), .wire_3_7_4_8_remainter(Remainder_out), .wire_3_06_07_curry(C_in), .wire_3_07_08_curry(C_out));
	div_cell cas_3_6 (.~wire_out_quotient_13(T_in), .divisor[6](Divisor_in), .wire_2_5_3_6_remainter(Remainder_in), .wire_3_6_4_7_remainter(Remainder_out), .wire_3_05_06_curry(C_in), .wire_3_06_07_curry(C_out));
	div_cell cas_3_5 (.~wire_out_quotient_13(T_in), .divisor[5](Divisor_in), .wire_2_4_3_5_remainter(Remainder_in), .wire_3_5_4_6_remainter(Remainder_out), .wire_3_04_05_curry(C_in), .wire_3_05_06_curry(C_out));
	div_cell cas_3_4 (.~wire_out_quotient_13(T_in), .divisor[4](Divisor_in), .wire_2_3_3_4_remainter(Remainder_in), .wire_3_4_4_5_remainter(Remainder_out), .wire_3_03_04_curry(C_in), .wire_3_04_05_curry(C_out));
	div_cell cas_3_3 (.~wire_out_quotient_13(T_in), .divisor[3](Divisor_in), .wire_2_2_3_3_remainter(Remainder_in), .wire_3_3_4_4_remainter(Remainder_out), .wire_3_02_03_curry(C_in), .wire_3_03_04_curry(C_out));
	div_cell cas_3_2 (.~wire_out_quotient_13(T_in), .divisor[2](Divisor_in), .wire_2_1_3_2_remainter(Remainder_in), .wire_3_2_4_3_remainter(Remainder_out), .wire_3_01_02_curry(C_in), .wire_3_02_03_curry(C_out));
	div_cell cas_3_1 (.~wire_out_quotient_13(T_in), .divisor[1](Divisor_in), .wire_2_0_3_1_remainter(Remainder_in), .wire_3_1_4_2_remainter(Remainder_out), .wire_3_00_01_curry(C_in), .wire_3_01_02_curry(C_out));

	div_cell cas_3_0 (.~wire_out_quotient_13(T_in), .divisor[0](Divisor_in), .dividend[13](Remainder_in), .wire_3_0_4_1_remainter(Remainder_out), .~wire_out_quotient_13(C_in), .wire_3_00_01_curry(C_out));

	//5th row
	div_cell cas_4_15 (.~wire_out_quotient_12(T_in), .divisor[15](Divisor_in), .wire_3_14_4_15_remainter(Remainder_in), .wire_out_quotient_11(Remainder_out), .wire_4_14_15_curry(C_in), .hang_4_wire_15(C_out));

	div_cell cas_4_14 (.~wire_out_quotient_12(T_in), .divisor[14](Divisor_in), .wire_3_13_4_14_remainter(Remainder_in), .wire_4_14_5_15_remainter(Remainder_out), .wire_4_13_14_curry(C_in), .wire_4_14_15_curry(C_out));
	div_cell cas_4_13 (.~wire_out_quotient_12(T_in), .divisor[13](Divisor_in), .wire_3_12_4_13_remainter(Remainder_in), .wire_4_13_5_14_remainter(Remainder_out), .wire_4_12_13_curry(C_in), .wire_4_13_14_curry(C_out));
	div_cell cas_4_12 (.~wire_out_quotient_12(T_in), .divisor[12](Divisor_in), .wire_3_11_4_12_remainter(Remainder_in), .wire_4_12_5_13_remainter(Remainder_out), .wire_4_11_12_curry(C_in), .wire_4_12_13_curry(C_out));
	div_cell cas_4_11 (.~wire_out_quotient_12(T_in), .divisor[11](Divisor_in), .wire_3_10_4_11_remainter(Remainder_in), .wire_4_11_5_12_remainter(Remainder_out), .wire_4_10_11_curry(C_in), .wire_4_11_12_curry(C_out));
	div_cell cas_4_10 (.~wire_out_quotient_12(T_in), .divisor[10](Divisor_in), .wire_3_9_4_10_remainter(Remainder_in), .wire_4_10_5_11_remainter(Remainder_out), .wire_4_09_10_curry(C_in), .wire_4_10_11_curry(C_out));
	div_cell cas_4_9 (.~wire_out_quotient_12(T_in), .divisor[9](Divisor_in), .wire_3_8_4_9_remainter(Remainder_in), .wire_4_9_5_10_remainter(Remainder_out), .wire_4_08_09_curry(C_in), .wire_4_09_10_curry(C_out));
	div_cell cas_4_8 (.~wire_out_quotient_12(T_in), .divisor[8](Divisor_in), .wire_3_7_4_8_remainter(Remainder_in), .wire_4_8_5_9_remainter(Remainder_out), .wire_4_07_08_curry(C_in), .wire_4_08_09_curry(C_out));
	div_cell cas_4_7 (.~wire_out_quotient_12(T_in), .divisor[7](Divisor_in), .wire_3_6_4_7_remainter(Remainder_in), .wire_4_7_5_8_remainter(Remainder_out), .wire_4_06_07_curry(C_in), .wire_4_07_08_curry(C_out));
	div_cell cas_4_6 (.~wire_out_quotient_12(T_in), .divisor[6](Divisor_in), .wire_3_5_4_6_remainter(Remainder_in), .wire_4_6_5_7_remainter(Remainder_out), .wire_4_05_06_curry(C_in), .wire_4_06_07_curry(C_out));
	div_cell cas_4_5 (.~wire_out_quotient_12(T_in), .divisor[5](Divisor_in), .wire_3_4_4_5_remainter(Remainder_in), .wire_4_5_5_6_remainter(Remainder_out), .wire_4_04_05_curry(C_in), .wire_4_05_06_curry(C_out));
	div_cell cas_4_4 (.~wire_out_quotient_12(T_in), .divisor[4](Divisor_in), .wire_3_3_4_4_remainter(Remainder_in), .wire_4_4_5_5_remainter(Remainder_out), .wire_4_03_04_curry(C_in), .wire_4_04_05_curry(C_out));
	div_cell cas_4_3 (.~wire_out_quotient_12(T_in), .divisor[3](Divisor_in), .wire_3_2_4_3_remainter(Remainder_in), .wire_4_3_5_4_remainter(Remainder_out), .wire_4_02_03_curry(C_in), .wire_4_03_04_curry(C_out));
	div_cell cas_4_2 (.~wire_out_quotient_12(T_in), .divisor[2](Divisor_in), .wire_3_1_4_2_remainter(Remainder_in), .wire_4_2_5_3_remainter(Remainder_out), .wire_4_01_02_curry(C_in), .wire_4_02_03_curry(C_out));
	div_cell cas_4_1 (.~wire_out_quotient_12(T_in), .divisor[1](Divisor_in), .wire_3_0_4_1_remainter(Remainder_in), .wire_4_1_5_2_remainter(Remainder_out), .wire_4_00_01_curry(C_in), .wire_4_01_02_curry(C_out));

	div_cell cas_4_0 (.~wire_out_quotient_12(T_in), .divisor[0](Divisor_in), .dividend[12](Remainder_in), .wire_4_0_5_1_remainter(Remainder_out), .~wire_out_quotient_12(C_in), .wire_4_00_01_curry(C_out));

	//6th row
	div_cell cas_5_15 (.~wire_out_quotient_11(T_in), .divisor[15](Divisor_in), .wire_4_14_5_15_remainter(Remainder_in), .wire_out_quotient_10(Remainder_out), .wire_5_14_15_curry(C_in), .hang_5_wire_15(C_out));

	div_cell cas_5_14 (.~wire_out_quotient_11(T_in), .divisor[14](Divisor_in), .wire_4_13_5_14_remainter(Remainder_in), .wire_5_14_6_15_remainter(Remainder_out), .wire_5_13_14_curry(C_in), .wire_5_14_15_curry(C_out));
	div_cell cas_5_13 (.~wire_out_quotient_11(T_in), .divisor[13](Divisor_in), .wire_4_12_5_13_remainter(Remainder_in), .wire_5_13_6_14_remainter(Remainder_out), .wire_5_12_13_curry(C_in), .wire_5_13_14_curry(C_out));
	div_cell cas_5_12 (.~wire_out_quotient_11(T_in), .divisor[12](Divisor_in), .wire_4_11_5_12_remainter(Remainder_in), .wire_5_12_6_13_remainter(Remainder_out), .wire_5_11_12_curry(C_in), .wire_5_12_13_curry(C_out));
	div_cell cas_5_11 (.~wire_out_quotient_11(T_in), .divisor[11](Divisor_in), .wire_4_10_5_11_remainter(Remainder_in), .wire_5_11_6_12_remainter(Remainder_out), .wire_5_10_11_curry(C_in), .wire_5_11_12_curry(C_out));
	div_cell cas_5_10 (.~wire_out_quotient_11(T_in), .divisor[10](Divisor_in), .wire_4_9_5_10_remainter(Remainder_in), .wire_5_10_6_11_remainter(Remainder_out), .wire_5_09_10_curry(C_in), .wire_5_10_11_curry(C_out));
	div_cell cas_5_9 (.~wire_out_quotient_11(T_in), .divisor[9](Divisor_in), .wire_4_8_5_9_remainter(Remainder_in), .wire_5_9_6_10_remainter(Remainder_out), .wire_5_08_09_curry(C_in), .wire_5_09_10_curry(C_out));
	div_cell cas_5_8 (.~wire_out_quotient_11(T_in), .divisor[8](Divisor_in), .wire_4_7_5_8_remainter(Remainder_in), .wire_5_8_6_9_remainter(Remainder_out), .wire_5_07_08_curry(C_in), .wire_5_08_09_curry(C_out));
	div_cell cas_5_7 (.~wire_out_quotient_11(T_in), .divisor[7](Divisor_in), .wire_4_6_5_7_remainter(Remainder_in), .wire_5_7_6_8_remainter(Remainder_out), .wire_5_06_07_curry(C_in), .wire_5_07_08_curry(C_out));
	div_cell cas_5_6 (.~wire_out_quotient_11(T_in), .divisor[6](Divisor_in), .wire_4_5_5_6_remainter(Remainder_in), .wire_5_6_6_7_remainter(Remainder_out), .wire_5_05_06_curry(C_in), .wire_5_06_07_curry(C_out));
	div_cell cas_5_5 (.~wire_out_quotient_11(T_in), .divisor[5](Divisor_in), .wire_4_4_5_5_remainter(Remainder_in), .wire_5_5_6_6_remainter(Remainder_out), .wire_5_04_05_curry(C_in), .wire_5_05_06_curry(C_out));
	div_cell cas_5_4 (.~wire_out_quotient_11(T_in), .divisor[4](Divisor_in), .wire_4_3_5_4_remainter(Remainder_in), .wire_5_4_6_5_remainter(Remainder_out), .wire_5_03_04_curry(C_in), .wire_5_04_05_curry(C_out));
	div_cell cas_5_3 (.~wire_out_quotient_11(T_in), .divisor[3](Divisor_in), .wire_4_2_5_3_remainter(Remainder_in), .wire_5_3_6_4_remainter(Remainder_out), .wire_5_02_03_curry(C_in), .wire_5_03_04_curry(C_out));
	div_cell cas_5_2 (.~wire_out_quotient_11(T_in), .divisor[2](Divisor_in), .wire_4_1_5_2_remainter(Remainder_in), .wire_5_2_6_3_remainter(Remainder_out), .wire_5_01_02_curry(C_in), .wire_5_02_03_curry(C_out));
	div_cell cas_5_1 (.~wire_out_quotient_11(T_in), .divisor[1](Divisor_in), .wire_4_0_5_1_remainter(Remainder_in), .wire_5_1_6_2_remainter(Remainder_out), .wire_5_00_01_curry(C_in), .wire_5_01_02_curry(C_out));

	div_cell cas_5_0 (.~wire_out_quotient_11(T_in), .divisor[0](Divisor_in), .dividend[11](Remainder_in), .wire_5_0_6_1_remainter(Remainder_out), .~wire_out_quotient_11(C_in), .wire_5_00_01_curry(C_out));

	//7th row
	div_cell cas_6_15 (.~wire_out_quotient_10(T_in), .divisor[15](Divisor_in), .wire_5_14_6_15_remainter(Remainder_in), .wire_out_quotient_9(Remainder_out), .wire_6_14_15_curry(C_in), .hang_6_wire_15(C_out));

	div_cell cas_6_14 (.~wire_out_quotient_10(T_in), .divisor[14](Divisor_in), .wire_5_13_6_14_remainter(Remainder_in), .wire_6_14_7_15_remainter(Remainder_out), .wire_6_13_14_curry(C_in), .wire_6_14_15_curry(C_out));
	div_cell cas_6_13 (.~wire_out_quotient_10(T_in), .divisor[13](Divisor_in), .wire_5_12_6_13_remainter(Remainder_in), .wire_6_13_7_14_remainter(Remainder_out), .wire_6_12_13_curry(C_in), .wire_6_13_14_curry(C_out));
	div_cell cas_6_12 (.~wire_out_quotient_10(T_in), .divisor[12](Divisor_in), .wire_5_11_6_12_remainter(Remainder_in), .wire_6_12_7_13_remainter(Remainder_out), .wire_6_11_12_curry(C_in), .wire_6_12_13_curry(C_out));
	div_cell cas_6_11 (.~wire_out_quotient_10(T_in), .divisor[11](Divisor_in), .wire_5_10_6_11_remainter(Remainder_in), .wire_6_11_7_12_remainter(Remainder_out), .wire_6_10_11_curry(C_in), .wire_6_11_12_curry(C_out));
	div_cell cas_6_10 (.~wire_out_quotient_10(T_in), .divisor[10](Divisor_in), .wire_5_9_6_10_remainter(Remainder_in), .wire_6_10_7_11_remainter(Remainder_out), .wire_6_09_10_curry(C_in), .wire_6_10_11_curry(C_out));
	div_cell cas_6_9 (.~wire_out_quotient_10(T_in), .divisor[9](Divisor_in), .wire_5_8_6_9_remainter(Remainder_in), .wire_6_9_7_10_remainter(Remainder_out), .wire_6_08_09_curry(C_in), .wire_6_09_10_curry(C_out));
	div_cell cas_6_8 (.~wire_out_quotient_10(T_in), .divisor[8](Divisor_in), .wire_5_7_6_8_remainter(Remainder_in), .wire_6_8_7_9_remainter(Remainder_out), .wire_6_07_08_curry(C_in), .wire_6_08_09_curry(C_out));
	div_cell cas_6_7 (.~wire_out_quotient_10(T_in), .divisor[7](Divisor_in), .wire_5_6_6_7_remainter(Remainder_in), .wire_6_7_7_8_remainter(Remainder_out), .wire_6_06_07_curry(C_in), .wire_6_07_08_curry(C_out));
	div_cell cas_6_6 (.~wire_out_quotient_10(T_in), .divisor[6](Divisor_in), .wire_5_5_6_6_remainter(Remainder_in), .wire_6_6_7_7_remainter(Remainder_out), .wire_6_05_06_curry(C_in), .wire_6_06_07_curry(C_out));
	div_cell cas_6_5 (.~wire_out_quotient_10(T_in), .divisor[5](Divisor_in), .wire_5_4_6_5_remainter(Remainder_in), .wire_6_5_7_6_remainter(Remainder_out), .wire_6_04_05_curry(C_in), .wire_6_05_06_curry(C_out));
	div_cell cas_6_4 (.~wire_out_quotient_10(T_in), .divisor[4](Divisor_in), .wire_5_3_6_4_remainter(Remainder_in), .wire_6_4_7_5_remainter(Remainder_out), .wire_6_03_04_curry(C_in), .wire_6_04_05_curry(C_out));
	div_cell cas_6_3 (.~wire_out_quotient_10(T_in), .divisor[3](Divisor_in), .wire_5_2_6_3_remainter(Remainder_in), .wire_6_3_7_4_remainter(Remainder_out), .wire_6_02_03_curry(C_in), .wire_6_03_04_curry(C_out));
	div_cell cas_6_2 (.~wire_out_quotient_10(T_in), .divisor[2](Divisor_in), .wire_5_1_6_2_remainter(Remainder_in), .wire_6_2_7_3_remainter(Remainder_out), .wire_6_01_02_curry(C_in), .wire_6_02_03_curry(C_out));
	div_cell cas_6_1 (.~wire_out_quotient_10(T_in), .divisor[1](Divisor_in), .wire_5_0_6_1_remainter(Remainder_in), .wire_6_1_7_2_remainter(Remainder_out), .wire_6_00_01_curry(C_in), .wire_6_01_02_curry(C_out));

	div_cell cas_6_0 (.~wire_out_quotient_10(T_in), .divisor[0](Divisor_in), .dividend[10](Remainder_in), .wire_6_0_7_1_remainter(Remainder_out), .~wire_out_quotient_10(C_in), .wire_6_00_01_curry(C_out));

	//8th row
	div_cell cas_7_15 (.~wire_out_quotient_9(T_in), .divisor[15](Divisor_in), .wire_6_14_7_15_remainter(Remainder_in), .wire_out_quotient_8(Remainder_out), .wire_7_14_15_curry(C_in), .hang_7_wire_15(C_out));

	div_cell cas_7_14 (.~wire_out_quotient_9(T_in), .divisor[14](Divisor_in), .wire_6_13_7_14_remainter(Remainder_in), .wire_7_14_8_15_remainter(Remainder_out), .wire_7_13_14_curry(C_in), .wire_7_14_15_curry(C_out));
	div_cell cas_7_13 (.~wire_out_quotient_9(T_in), .divisor[13](Divisor_in), .wire_6_12_7_13_remainter(Remainder_in), .wire_7_13_8_14_remainter(Remainder_out), .wire_7_12_13_curry(C_in), .wire_7_13_14_curry(C_out));
	div_cell cas_7_12 (.~wire_out_quotient_9(T_in), .divisor[12](Divisor_in), .wire_6_11_7_12_remainter(Remainder_in), .wire_7_12_8_13_remainter(Remainder_out), .wire_7_11_12_curry(C_in), .wire_7_12_13_curry(C_out));
	div_cell cas_7_11 (.~wire_out_quotient_9(T_in), .divisor[11](Divisor_in), .wire_6_10_7_11_remainter(Remainder_in), .wire_7_11_8_12_remainter(Remainder_out), .wire_7_10_11_curry(C_in), .wire_7_11_12_curry(C_out));
	div_cell cas_7_10 (.~wire_out_quotient_9(T_in), .divisor[10](Divisor_in), .wire_6_9_7_10_remainter(Remainder_in), .wire_7_10_8_11_remainter(Remainder_out), .wire_7_09_10_curry(C_in), .wire_7_10_11_curry(C_out));
	div_cell cas_7_9 (.~wire_out_quotient_9(T_in), .divisor[9](Divisor_in), .wire_6_8_7_9_remainter(Remainder_in), .wire_7_9_8_10_remainter(Remainder_out), .wire_7_08_09_curry(C_in), .wire_7_09_10_curry(C_out));
	div_cell cas_7_8 (.~wire_out_quotient_9(T_in), .divisor[8](Divisor_in), .wire_6_7_7_8_remainter(Remainder_in), .wire_7_8_8_9_remainter(Remainder_out), .wire_7_07_08_curry(C_in), .wire_7_08_09_curry(C_out));
	div_cell cas_7_7 (.~wire_out_quotient_9(T_in), .divisor[7](Divisor_in), .wire_6_6_7_7_remainter(Remainder_in), .wire_7_7_8_8_remainter(Remainder_out), .wire_7_06_07_curry(C_in), .wire_7_07_08_curry(C_out));
	div_cell cas_7_6 (.~wire_out_quotient_9(T_in), .divisor[6](Divisor_in), .wire_6_5_7_6_remainter(Remainder_in), .wire_7_6_8_7_remainter(Remainder_out), .wire_7_05_06_curry(C_in), .wire_7_06_07_curry(C_out));
	div_cell cas_7_5 (.~wire_out_quotient_9(T_in), .divisor[5](Divisor_in), .wire_6_4_7_5_remainter(Remainder_in), .wire_7_5_8_6_remainter(Remainder_out), .wire_7_04_05_curry(C_in), .wire_7_05_06_curry(C_out));
	div_cell cas_7_4 (.~wire_out_quotient_9(T_in), .divisor[4](Divisor_in), .wire_6_3_7_4_remainter(Remainder_in), .wire_7_4_8_5_remainter(Remainder_out), .wire_7_03_04_curry(C_in), .wire_7_04_05_curry(C_out));
	div_cell cas_7_3 (.~wire_out_quotient_9(T_in), .divisor[3](Divisor_in), .wire_6_2_7_3_remainter(Remainder_in), .wire_7_3_8_4_remainter(Remainder_out), .wire_7_02_03_curry(C_in), .wire_7_03_04_curry(C_out));
	div_cell cas_7_2 (.~wire_out_quotient_9(T_in), .divisor[2](Divisor_in), .wire_6_1_7_2_remainter(Remainder_in), .wire_7_2_8_3_remainter(Remainder_out), .wire_7_01_02_curry(C_in), .wire_7_02_03_curry(C_out));
	div_cell cas_7_1 (.~wire_out_quotient_9(T_in), .divisor[1](Divisor_in), .wire_6_0_7_1_remainter(Remainder_in), .wire_7_1_8_2_remainter(Remainder_out), .wire_7_00_01_curry(C_in), .wire_7_01_02_curry(C_out));
	
	div_cell cas_7_0 (.~wire_out_quotient_9(T_in), .divisor[0](Divisor_in), .dividend[9](Remainder_in), .wire_7_0_8_1_remainter(Remainder_out), .~wire_out_quotient_9(C_in), .wire_7_00_01_curry(C_out));

	//9th row
	div_cell cas_8_15 (.~wire_out_quotient_8(T_in), .divisor[15](Divisor_in), .wire_7_14_8_15_remainter(Remainder_in), .wire_out_quotient_7(Remainder_out), .wire_8_14_15_curry(C_in), .hang_8_wire_15(C_out));

	div_cell cas_8_14 (.~wire_out_quotient_8(T_in), .divisor[14](Divisor_in), .wire_7_13_8_14_remainter(Remainder_in), .wire_8_14_9_15_remainter(Remainder_out), .wire_8_13_14_curry(C_in), .wire_8_14_15_curry(C_out));
	div_cell cas_8_13 (.~wire_out_quotient_8(T_in), .divisor[13](Divisor_in), .wire_7_12_8_13_remainter(Remainder_in), .wire_8_13_9_14_remainter(Remainder_out), .wire_8_12_13_curry(C_in), .wire_8_13_14_curry(C_out));
	div_cell cas_8_12 (.~wire_out_quotient_8(T_in), .divisor[12](Divisor_in), .wire_7_11_8_12_remainter(Remainder_in), .wire_8_12_9_13_remainter(Remainder_out), .wire_8_11_12_curry(C_in), .wire_8_12_13_curry(C_out));
	div_cell cas_8_11 (.~wire_out_quotient_8(T_in), .divisor[11](Divisor_in), .wire_7_10_8_11_remainter(Remainder_in), .wire_8_11_9_12_remainter(Remainder_out), .wire_8_10_11_curry(C_in), .wire_8_11_12_curry(C_out));
	div_cell cas_8_10 (.~wire_out_quotient_8(T_in), .divisor[10](Divisor_in), .wire_7_9_8_10_remainter(Remainder_in), .wire_8_10_9_11_remainter(Remainder_out), .wire_8_09_10_curry(C_in), .wire_8_10_11_curry(C_out));
	div_cell cas_8_9 (.~wire_out_quotient_8(T_in), .divisor[9](Divisor_in), .wire_7_8_8_9_remainter(Remainder_in), .wire_8_9_9_10_remainter(Remainder_out), .wire_8_08_09_curry(C_in), .wire_8_09_10_curry(C_out));
	div_cell cas_8_8 (.~wire_out_quotient_8(T_in), .divisor[8](Divisor_in), .wire_7_7_8_8_remainter(Remainder_in), .wire_8_8_9_9_remainter(Remainder_out), .wire_8_07_08_curry(C_in), .wire_8_08_09_curry(C_out));
	div_cell cas_8_7 (.~wire_out_quotient_8(T_in), .divisor[7](Divisor_in), .wire_7_6_8_7_remainter(Remainder_in), .wire_8_7_9_8_remainter(Remainder_out), .wire_8_06_07_curry(C_in), .wire_8_07_08_curry(C_out));
	div_cell cas_8_6 (.~wire_out_quotient_8(T_in), .divisor[6](Divisor_in), .wire_7_5_8_6_remainter(Remainder_in), .wire_8_6_9_7_remainter(Remainder_out), .wire_8_05_06_curry(C_in), .wire_8_06_07_curry(C_out));
	div_cell cas_8_5 (.~wire_out_quotient_8(T_in), .divisor[5](Divisor_in), .wire_7_4_8_5_remainter(Remainder_in), .wire_8_5_9_6_remainter(Remainder_out), .wire_8_04_05_curry(C_in), .wire_8_05_06_curry(C_out));
	div_cell cas_8_4 (.~wire_out_quotient_8(T_in), .divisor[4](Divisor_in), .wire_7_3_8_4_remainter(Remainder_in), .wire_8_4_9_5_remainter(Remainder_out), .wire_8_03_04_curry(C_in), .wire_8_04_05_curry(C_out));
	div_cell cas_8_3 (.~wire_out_quotient_8(T_in), .divisor[3](Divisor_in), .wire_7_2_8_3_remainter(Remainder_in), .wire_8_3_9_4_remainter(Remainder_out), .wire_8_02_03_curry(C_in), .wire_8_03_04_curry(C_out));
	div_cell cas_8_2 (.~wire_out_quotient_8(T_in), .divisor[2](Divisor_in), .wire_7_1_8_2_remainter(Remainder_in), .wire_8_2_9_3_remainter(Remainder_out), .wire_8_01_02_curry(C_in), .wire_8_02_03_curry(C_out));
	div_cell cas_8_1 (.~wire_out_quotient_8(T_in), .divisor[1](Divisor_in), .wire_7_0_8_1_remainter(Remainder_in), .wire_8_1_9_2_remainter(Remainder_out), .wire_8_00_01_curry(C_in), .wire_8_01_02_curry(C_out));
	
	div_cell cas_8_0 (.~wire_out_quotient_8(T_in), .divisor[0](Divisor_in), .dividend[8](Remainder_in), .wire_8_0_9_1_remainter(Remainder_out), .~wire_out_quotient_8(C_in), .wire_8_00_01_curry(C_out));

	//10th row
	div_cell cas_9_15 (.~wire_out_quotient_7(T_in), .divisor[15](Divisor_in), .wire_8_14_9_15_remainter(Remainder_in), .wire_out_quotient_6(Remainder_out), .wire_9_14_15_curry(C_in), .hang_9_wire_15(C_out));

	div_cell cas_9_14 (.~wire_out_quotient_7(T_in), .divisor[14](Divisor_in), .wire_8_13_9_14_remainter(Remainder_in), .wire_9_14_10_15_remainter(Remainder_out), .wire_9_13_14_curry(C_in), .wire_9_14_15_curry(C_out));
	div_cell cas_9_13 (.~wire_out_quotient_7(T_in), .divisor[13](Divisor_in), .wire_8_12_9_13_remainter(Remainder_in), .wire_9_13_10_14_remainter(Remainder_out), .wire_9_12_13_curry(C_in), .wire_9_13_14_curry(C_out));
	div_cell cas_9_12 (.~wire_out_quotient_7(T_in), .divisor[12](Divisor_in), .wire_8_11_9_12_remainter(Remainder_in), .wire_9_12_10_13_remainter(Remainder_out), .wire_9_11_12_curry(C_in), .wire_9_12_13_curry(C_out));
	div_cell cas_9_11 (.~wire_out_quotient_7(T_in), .divisor[11](Divisor_in), .wire_8_10_9_11_remainter(Remainder_in), .wire_9_11_10_12_remainter(Remainder_out), .wire_9_10_11_curry(C_in), .wire_9_11_12_curry(C_out));
	div_cell cas_9_10 (.~wire_out_quotient_7(T_in), .divisor[10](Divisor_in), .wire_8_9_9_10_remainter(Remainder_in), .wire_9_10_10_11_remainter(Remainder_out), .wire_9_09_10_curry(C_in), .wire_9_10_11_curry(C_out));
	div_cell cas_9_9 (.~wire_out_quotient_7(T_in), .divisor[9](Divisor_in), .wire_8_8_9_9_remainter(Remainder_in), .wire_9_9_10_10_remainter(Remainder_out), .wire_9_08_09_curry(C_in), .wire_9_09_10_curry(C_out));
	div_cell cas_9_8 (.~wire_out_quotient_7(T_in), .divisor[8](Divisor_in), .wire_8_7_9_8_remainter(Remainder_in), .wire_9_8_10_9_remainter(Remainder_out), .wire_9_07_08_curry(C_in), .wire_9_08_09_curry(C_out));
	div_cell cas_9_7 (.~wire_out_quotient_7(T_in), .divisor[7](Divisor_in), .wire_8_6_9_7_remainter(Remainder_in), .wire_9_7_10_8_remainter(Remainder_out), .wire_9_06_07_curry(C_in), .wire_9_07_08_curry(C_out));
	div_cell cas_9_6 (.~wire_out_quotient_7(T_in), .divisor[6](Divisor_in), .wire_8_5_9_6_remainter(Remainder_in), .wire_9_6_10_7_remainter(Remainder_out), .wire_9_05_06_curry(C_in), .wire_9_06_07_curry(C_out));
	div_cell cas_9_5 (.~wire_out_quotient_7(T_in), .divisor[5](Divisor_in), .wire_8_4_9_5_remainter(Remainder_in), .wire_9_5_10_6_remainter(Remainder_out), .wire_9_04_05_curry(C_in), .wire_9_05_06_curry(C_out));
	div_cell cas_9_4 (.~wire_out_quotient_7(T_in), .divisor[4](Divisor_in), .wire_8_3_9_4_remainter(Remainder_in), .wire_9_4_10_5_remainter(Remainder_out), .wire_9_03_04_curry(C_in), .wire_9_04_05_curry(C_out));
	div_cell cas_9_3 (.~wire_out_quotient_7(T_in), .divisor[3](Divisor_in), .wire_8_2_9_3_remainter(Remainder_in), .wire_9_3_10_4_remainter(Remainder_out), .wire_9_02_03_curry(C_in), .wire_9_03_04_curry(C_out));
	div_cell cas_9_2 (.~wire_out_quotient_7(T_in), .divisor[2](Divisor_in), .wire_8_1_9_2_remainter(Remainder_in), .wire_9_2_10_3_remainter(Remainder_out), .wire_9_01_02_curry(C_in), .wire_9_02_03_curry(C_out));
	div_cell cas_9_1 (.~wire_out_quotient_7(T_in), .divisor[1](Divisor_in), .wire_8_0_9_1_remainter(Remainder_in), .wire_9_1_10_2_remainter(Remainder_out), .wire_9_00_01_curry(C_in), .wire_9_01_02_curry(C_out));
	
	div_cell cas_9_0 (.~wire_out_quotient_7(T_in), .divisor[0](Divisor_in), .dividend[7](Remainder_in), .wire_9_0_10_1_remainter(Remainder_out), .~wire_out_quotient_7(C_in), .wire_9_00_01_curry(C_out));

	//11th row
	div_cell cas_10_15 (.~wire_out_quotient_6(T_in), .divisor[15](Divisor_in), .wire_9_14_10_15_remainter(Remainder_in), .wire_out_quotient_5(Remainder_out), .wire_10_14_15_curry(C_in), .hang_10_wire_15(C_out));

	div_cell cas_10_14 (.~wire_out_quotient_6(T_in), .divisor[14](Divisor_in), .wire_9_13_10_14_remainter(Remainder_in), .wire_10_14_11_15_remainter(Remainder_out), .wire_10_13_14_curry(C_in), .wire_10_14_15_curry(C_out));
	div_cell cas_10_13 (.~wire_out_quotient_6(T_in), .divisor[13](Divisor_in), .wire_9_12_10_13_remainter(Remainder_in), .wire_10_13_11_14_remainter(Remainder_out), .wire_10_12_13_curry(C_in), .wire_10_13_14_curry(C_out));
	div_cell cas_10_12 (.~wire_out_quotient_6(T_in), .divisor[12](Divisor_in), .wire_9_11_10_12_remainter(Remainder_in), .wire_10_12_11_13_remainter(Remainder_out), .wire_10_11_12_curry(C_in), .wire_10_12_13_curry(C_out));
	div_cell cas_10_11 (.~wire_out_quotient_6(T_in), .divisor[11](Divisor_in), .wire_9_10_10_11_remainter(Remainder_in), .wire_10_11_11_12_remainter(Remainder_out), .wire_10_10_11_curry(C_in), .wire_10_11_12_curry(C_out));
	div_cell cas_10_10 (.~wire_out_quotient_6(T_in), .divisor[10](Divisor_in), .wire_9_9_10_10_remainter(Remainder_in), .wire_10_10_11_11_remainter(Remainder_out), .wire_10_09_10_curry(C_in), .wire_10_10_11_curry(C_out));
	div_cell cas_10_9 (.~wire_out_quotient_6(T_in), .divisor[9](Divisor_in), .wire_9_8_10_9_remainter(Remainder_in), .wire_10_9_11_10_remainter(Remainder_out), .wire_10_08_09_curry(C_in), .wire_10_09_10_curry(C_out));
	div_cell cas_10_8 (.~wire_out_quotient_6(T_in), .divisor[8](Divisor_in), .wire_9_7_10_8_remainter(Remainder_in), .wire_10_8_11_9_remainter(Remainder_out), .wire_10_07_08_curry(C_in), .wire_10_08_09_curry(C_out));
	div_cell cas_10_7 (.~wire_out_quotient_6(T_in), .divisor[7](Divisor_in), .wire_9_6_10_7_remainter(Remainder_in), .wire_10_7_11_8_remainter(Remainder_out), .wire_10_06_07_curry(C_in), .wire_10_07_08_curry(C_out));
	div_cell cas_10_6 (.~wire_out_quotient_6(T_in), .divisor[6](Divisor_in), .wire_9_5_10_6_remainter(Remainder_in), .wire_10_6_11_7_remainter(Remainder_out), .wire_10_05_06_curry(C_in), .wire_10_06_07_curry(C_out));
	div_cell cas_10_5 (.~wire_out_quotient_6(T_in), .divisor[5](Divisor_in), .wire_9_4_10_5_remainter(Remainder_in), .wire_10_5_11_6_remainter(Remainder_out), .wire_10_04_05_curry(C_in), .wire_10_05_06_curry(C_out));
	div_cell cas_10_4 (.~wire_out_quotient_6(T_in), .divisor[4](Divisor_in), .wire_9_3_10_4_remainter(Remainder_in), .wire_10_4_11_5_remainter(Remainder_out), .wire_10_03_04_curry(C_in), .wire_10_04_05_curry(C_out));
	div_cell cas_10_3 (.~wire_out_quotient_6(T_in), .divisor[3](Divisor_in), .wire_9_2_10_3_remainter(Remainder_in), .wire_10_3_11_4_remainter(Remainder_out), .wire_10_02_03_curry(C_in), .wire_10_03_04_curry(C_out));
	div_cell cas_10_2 (.~wire_out_quotient_6(T_in), .divisor[2](Divisor_in), .wire_9_1_10_2_remainter(Remainder_in), .wire_10_2_11_3_remainter(Remainder_out), .wire_10_01_02_curry(C_in), .wire_10_02_03_curry(C_out));
	div_cell cas_10_1 (.~wire_out_quotient_6(T_in), .divisor[1](Divisor_in), .wire_9_0_10_1_remainter(Remainder_in), .wire_10_1_11_2_remainter(Remainder_out), .wire_10_00_01_curry(C_in), .wire_10_01_02_curry(C_out));
	
	div_cell cas_10_0 (.~wire_out_quotient_6(T_in), .divisor[0](Divisor_in), .dividend[6](Remainder_in), .wire_10_0_11_1_remainter(Remainder_out), .~wire_out_quotient_6(C_in), .wire_10_00_01_curry(C_out));

	//12th row
	div_cell cas_11_15 (.~wire_out_quotient_5(T_in), .divisor[15](Divisor_in), .wire_10_14_11_15_remainter(Remainder_in), .wire_out_quotient_4(Remainder_out), .wire_11_14_15_curry(C_in), .hang_11_wire_15(C_out));

	div_cell cas_11_14 (.~wire_out_quotient_5(T_in), .divisor[14](Divisor_in), .wire_10_13_11_14_remainter(Remainder_in), .wire_11_14_12_15_remainter(Remainder_out), .wire_11_13_14_curry(C_in), .wire_11_14_15_curry(C_out));
	div_cell cas_11_13 (.~wire_out_quotient_5(T_in), .divisor[13](Divisor_in), .wire_10_12_11_13_remainter(Remainder_in), .wire_11_13_12_14_remainter(Remainder_out), .wire_11_12_13_curry(C_in), .wire_11_13_14_curry(C_out));
	div_cell cas_11_12 (.~wire_out_quotient_5(T_in), .divisor[12](Divisor_in), .wire_10_11_11_12_remainter(Remainder_in), .wire_11_12_12_13_remainter(Remainder_out), .wire_11_11_12_curry(C_in), .wire_11_12_13_curry(C_out));
	div_cell cas_11_11 (.~wire_out_quotient_5(T_in), .divisor[11](Divisor_in), .wire_10_10_11_11_remainter(Remainder_in), .wire_11_11_12_12_remainter(Remainder_out), .wire_11_10_11_curry(C_in), .wire_11_11_12_curry(C_out));
	div_cell cas_11_10 (.~wire_out_quotient_5(T_in), .divisor[10](Divisor_in), .wire_10_9_11_10_remainter(Remainder_in), .wire_11_10_12_11_remainter(Remainder_out), .wire_11_09_10_curry(C_in), .wire_11_10_11_curry(C_out));
	div_cell cas_11_9 (.~wire_out_quotient_5(T_in), .divisor[9](Divisor_in), .wire_10_8_11_9_remainter(Remainder_in), .wire_11_9_12_10_remainter(Remainder_out), .wire_11_08_09_curry(C_in), .wire_11_09_10_curry(C_out));
	div_cell cas_11_8 (.~wire_out_quotient_5(T_in), .divisor[8](Divisor_in), .wire_10_7_11_8_remainter(Remainder_in), .wire_11_8_12_9_remainter(Remainder_out), .wire_11_07_08_curry(C_in), .wire_11_08_09_curry(C_out));
	div_cell cas_11_7 (.~wire_out_quotient_5(T_in), .divisor[7](Divisor_in), .wire_10_6_11_7_remainter(Remainder_in), .wire_11_7_12_8_remainter(Remainder_out), .wire_11_06_07_curry(C_in), .wire_11_07_08_curry(C_out));
	div_cell cas_11_6 (.~wire_out_quotient_5(T_in), .divisor[6](Divisor_in), .wire_10_5_11_6_remainter(Remainder_in), .wire_11_6_12_7_remainter(Remainder_out), .wire_11_05_06_curry(C_in), .wire_11_06_07_curry(C_out));
	div_cell cas_11_5 (.~wire_out_quotient_5(T_in), .divisor[5](Divisor_in), .wire_10_4_11_5_remainter(Remainder_in), .wire_11_5_12_6_remainter(Remainder_out), .wire_11_04_05_curry(C_in), .wire_11_05_06_curry(C_out));
	div_cell cas_11_4 (.~wire_out_quotient_5(T_in), .divisor[4](Divisor_in), .wire_10_3_11_4_remainter(Remainder_in), .wire_11_4_12_5_remainter(Remainder_out), .wire_11_03_04_curry(C_in), .wire_11_04_05_curry(C_out));
	div_cell cas_11_3 (.~wire_out_quotient_5(T_in), .divisor[3](Divisor_in), .wire_10_2_11_3_remainter(Remainder_in), .wire_11_3_12_4_remainter(Remainder_out), .wire_11_02_03_curry(C_in), .wire_11_03_04_curry(C_out));
	div_cell cas_11_2 (.~wire_out_quotient_5(T_in), .divisor[2](Divisor_in), .wire_10_1_11_2_remainter(Remainder_in), .wire_11_2_12_3_remainter(Remainder_out), .wire_11_01_02_curry(C_in), .wire_11_02_03_curry(C_out));
	div_cell cas_11_1 (.~wire_out_quotient_5(T_in), .divisor[1](Divisor_in), .wire_10_0_11_1_remainter(Remainder_in), .wire_11_1_12_2_remainter(Remainder_out), .wire_11_00_01_curry(C_in), .wire_11_01_02_curry(C_out));
	
	div_cell cas_11_0 (.~wire_out_quotient_5(T_in), .divisor[0](Divisor_in), .dividend[5](Remainder_in), .wire_11_0_12_1_remainter(Remainder_out), .~wire_out_quotient_5(C_in), .wire_11_00_01_curry(C_out));

	//13th row
	div_cell cas_12_15 (.~wire_out_quotient_4(T_in), .divisor[15](Divisor_in), .wire_11_14_12_15_remainter(Remainder_in), .wire_out_quotient_3(Remainder_out), .wire_12_14_15_curry(C_in), .hang_12_wire_15(C_out));

	div_cell cas_12_14 (.~wire_out_quotient_4(T_in), .divisor[14](Divisor_in), .wire_11_13_12_14_remainter(Remainder_in), .wire_12_14_13_15_remainter(Remainder_out), .wire_12_13_14_curry(C_in), .wire_12_14_15_curry(C_out));
	div_cell cas_12_13 (.~wire_out_quotient_4(T_in), .divisor[13](Divisor_in), .wire_11_12_12_13_remainter(Remainder_in), .wire_12_13_13_14_remainter(Remainder_out), .wire_12_12_13_curry(C_in), .wire_12_13_14_curry(C_out));
	div_cell cas_12_12 (.~wire_out_quotient_4(T_in), .divisor[12](Divisor_in), .wire_11_11_12_12_remainter(Remainder_in), .wire_12_12_13_13_remainter(Remainder_out), .wire_12_11_12_curry(C_in), .wire_12_12_13_curry(C_out));
	div_cell cas_12_11 (.~wire_out_quotient_4(T_in), .divisor[11](Divisor_in), .wire_11_10_12_11_remainter(Remainder_in), .wire_12_11_13_12_remainter(Remainder_out), .wire_12_10_11_curry(C_in), .wire_12_11_12_curry(C_out));
	div_cell cas_12_10 (.~wire_out_quotient_4(T_in), .divisor[10](Divisor_in), .wire_11_9_12_10_remainter(Remainder_in), .wire_12_10_13_11_remainter(Remainder_out), .wire_12_09_10_curry(C_in), .wire_12_10_11_curry(C_out));
	div_cell cas_12_9 (.~wire_out_quotient_4(T_in), .divisor[9](Divisor_in), .wire_11_8_12_9_remainter(Remainder_in), .wire_12_9_13_10_remainter(Remainder_out), .wire_12_08_09_curry(C_in), .wire_12_09_10_curry(C_out));
	div_cell cas_12_8 (.~wire_out_quotient_4(T_in), .divisor[8](Divisor_in), .wire_11_7_12_8_remainter(Remainder_in), .wire_12_8_13_9_remainter(Remainder_out), .wire_12_07_08_curry(C_in), .wire_12_08_09_curry(C_out));
	div_cell cas_12_7 (.~wire_out_quotient_4(T_in), .divisor[7](Divisor_in), .wire_11_6_12_7_remainter(Remainder_in), .wire_12_7_13_8_remainter(Remainder_out), .wire_12_06_07_curry(C_in), .wire_12_07_08_curry(C_out));
	div_cell cas_12_6 (.~wire_out_quotient_4(T_in), .divisor[6](Divisor_in), .wire_11_5_12_6_remainter(Remainder_in), .wire_12_6_13_7_remainter(Remainder_out), .wire_12_05_06_curry(C_in), .wire_12_06_07_curry(C_out));
	div_cell cas_12_5 (.~wire_out_quotient_4(T_in), .divisor[5](Divisor_in), .wire_11_4_12_5_remainter(Remainder_in), .wire_12_5_13_6_remainter(Remainder_out), .wire_12_04_05_curry(C_in), .wire_12_05_06_curry(C_out));
	div_cell cas_12_4 (.~wire_out_quotient_4(T_in), .divisor[4](Divisor_in), .wire_11_3_12_4_remainter(Remainder_in), .wire_12_4_13_5_remainter(Remainder_out), .wire_12_03_04_curry(C_in), .wire_12_04_05_curry(C_out));
	div_cell cas_12_3 (.~wire_out_quotient_4(T_in), .divisor[3](Divisor_in), .wire_11_2_12_3_remainter(Remainder_in), .wire_12_3_13_4_remainter(Remainder_out), .wire_12_02_03_curry(C_in), .wire_12_03_04_curry(C_out));
	div_cell cas_12_2 (.~wire_out_quotient_4(T_in), .divisor[2](Divisor_in), .wire_11_1_12_2_remainter(Remainder_in), .wire_12_2_13_3_remainter(Remainder_out), .wire_12_01_02_curry(C_in), .wire_12_02_03_curry(C_out));
	div_cell cas_12_1 (.~wire_out_quotient_4(T_in), .divisor[1](Divisor_in), .wire_11_0_12_1_remainter(Remainder_in), .wire_12_1_13_2_remainter(Remainder_out), .wire_12_00_01_curry(C_in), .wire_12_01_02_curry(C_out));
	
	div_cell cas_12_0 (.~wire_out_quotient_4(T_in), .divisor[0](Divisor_in), .dividend[4](Remainder_in), .wire_12_0_13_1_remainter(Remainder_out), .~wire_out_quotient_4(C_in), .wire_12_00_01_curry(C_out));

	//14th row
	div_cell cas_13_15 (.~wire_out_quotient_3(T_in), .divisor[15](Divisor_in), .wire_12_14_13_15_remainter(Remainder_in), .wire_out_quotient_2(Remainder_out), .wire_13_14_15_curry(C_in), .hang_13_wire_15(C_out));

	div_cell cas_13_14 (.~wire_out_quotient_3(T_in), .divisor[14](Divisor_in), .wire_12_13_13_14_remainter(Remainder_in), .wire_13_14_14_15_remainter(Remainder_out), .wire_13_13_14_curry(C_in), .wire_13_14_15_curry(C_out));
	div_cell cas_13_13 (.~wire_out_quotient_3(T_in), .divisor[13](Divisor_in), .wire_12_12_13_13_remainter(Remainder_in), .wire_13_13_14_14_remainter(Remainder_out), .wire_13_12_13_curry(C_in), .wire_13_13_14_curry(C_out));
	div_cell cas_13_12 (.~wire_out_quotient_3(T_in), .divisor[12](Divisor_in), .wire_12_11_13_12_remainter(Remainder_in), .wire_13_12_14_13_remainter(Remainder_out), .wire_13_11_12_curry(C_in), .wire_13_12_13_curry(C_out));
	div_cell cas_13_11 (.~wire_out_quotient_3(T_in), .divisor[11](Divisor_in), .wire_12_10_13_11_remainter(Remainder_in), .wire_13_11_14_12_remainter(Remainder_out), .wire_13_10_11_curry(C_in), .wire_13_11_12_curry(C_out));
	div_cell cas_13_10 (.~wire_out_quotient_3(T_in), .divisor[10](Divisor_in), .wire_12_9_13_10_remainter(Remainder_in), .wire_13_10_14_11_remainter(Remainder_out), .wire_13_09_10_curry(C_in), .wire_13_10_11_curry(C_out));
	div_cell cas_13_9 (.~wire_out_quotient_3(T_in), .divisor[9](Divisor_in), .wire_12_8_13_9_remainter(Remainder_in), .wire_13_9_14_10_remainter(Remainder_out), .wire_13_08_09_curry(C_in), .wire_13_09_10_curry(C_out));
	div_cell cas_13_8 (.~wire_out_quotient_3(T_in), .divisor[8](Divisor_in), .wire_12_7_13_8_remainter(Remainder_in), .wire_13_8_14_9_remainter(Remainder_out), .wire_13_07_08_curry(C_in), .wire_13_08_09_curry(C_out));
	div_cell cas_13_7 (.~wire_out_quotient_3(T_in), .divisor[7](Divisor_in), .wire_12_6_13_7_remainter(Remainder_in), .wire_13_7_14_8_remainter(Remainder_out), .wire_13_06_07_curry(C_in), .wire_13_07_08_curry(C_out));
	div_cell cas_13_6 (.~wire_out_quotient_3(T_in), .divisor[6](Divisor_in), .wire_12_5_13_6_remainter(Remainder_in), .wire_13_6_14_7_remainter(Remainder_out), .wire_13_05_06_curry(C_in), .wire_13_06_07_curry(C_out));
	div_cell cas_13_5 (.~wire_out_quotient_3(T_in), .divisor[5](Divisor_in), .wire_12_4_13_5_remainter(Remainder_in), .wire_13_5_14_6_remainter(Remainder_out), .wire_13_04_05_curry(C_in), .wire_13_05_06_curry(C_out));
	div_cell cas_13_4 (.~wire_out_quotient_3(T_in), .divisor[4](Divisor_in), .wire_12_3_13_4_remainter(Remainder_in), .wire_13_4_14_5_remainter(Remainder_out), .wire_13_03_04_curry(C_in), .wire_13_04_05_curry(C_out));
	div_cell cas_13_3 (.~wire_out_quotient_3(T_in), .divisor[3](Divisor_in), .wire_12_2_13_3_remainter(Remainder_in), .wire_13_3_14_4_remainter(Remainder_out), .wire_13_02_03_curry(C_in), .wire_13_03_04_curry(C_out));
	div_cell cas_13_2 (.~wire_out_quotient_3(T_in), .divisor[2](Divisor_in), .wire_12_1_13_2_remainter(Remainder_in), .wire_13_2_14_3_remainter(Remainder_out), .wire_13_01_02_curry(C_in), .wire_13_02_03_curry(C_out));
	div_cell cas_13_1 (.~wire_out_quotient_3(T_in), .divisor[1](Divisor_in), .wire_12_0_13_1_remainter(Remainder_in), .wire_13_1_14_2_remainter(Remainder_out), .wire_13_00_01_curry(C_in), .wire_13_01_02_curry(C_out));
	
	div_cell cas_13_0 (.~wire_out_quotient_3(T_in), .divisor[0](Divisor_in), .dividend[3](Remainder_in), .wire_13_0_14_1_remainter(Remainder_out), .~wire_out_quotient_3(C_in), .wire_13_00_01_curry(C_out));

	//15th row
	div_cell cas_13_15 (.~wire_out_quotient_3(T_in), .divisor[15](Divisor_in), .wire_12_14_13_15_remainter(Remainder_in), .wire_out_quotient_2(Remainder_out), .wire_13_14_15_curry(C_in), .hang_13_wire_15(C_out));

	div_cell cas_13_14 (.~wire_out_quotient_3(T_in), .divisor[14](Divisor_in), .wire_12_13_13_14_remainter(Remainder_in), .wire_13_14_14_15_remainter(Remainder_out), .wire_13_13_14_curry(C_in), .wire_13_14_15_curry(C_out));
	div_cell cas_13_13 (.~wire_out_quotient_3(T_in), .divisor[13](Divisor_in), .wire_12_12_13_13_remainter(Remainder_in), .wire_13_13_14_14_remainter(Remainder_out), .wire_13_12_13_curry(C_in), .wire_13_13_14_curry(C_out));
	div_cell cas_13_12 (.~wire_out_quotient_3(T_in), .divisor[12](Divisor_in), .wire_12_11_13_12_remainter(Remainder_in), .wire_13_12_14_13_remainter(Remainder_out), .wire_13_11_12_curry(C_in), .wire_13_12_13_curry(C_out));
	div_cell cas_13_11 (.~wire_out_quotient_3(T_in), .divisor[11](Divisor_in), .wire_12_10_13_11_remainter(Remainder_in), .wire_13_11_14_12_remainter(Remainder_out), .wire_13_10_11_curry(C_in), .wire_13_11_12_curry(C_out));
	div_cell cas_13_10 (.~wire_out_quotient_3(T_in), .divisor[10](Divisor_in), .wire_12_9_13_10_remainter(Remainder_in), .wire_13_10_14_11_remainter(Remainder_out), .wire_13_09_10_curry(C_in), .wire_13_10_11_curry(C_out));
	div_cell cas_13_9 (.~wire_out_quotient_3(T_in), .divisor[9](Divisor_in), .wire_12_8_13_9_remainter(Remainder_in), .wire_13_9_14_10_remainter(Remainder_out), .wire_13_08_09_curry(C_in), .wire_13_09_10_curry(C_out));
	div_cell cas_13_8 (.~wire_out_quotient_3(T_in), .divisor[8](Divisor_in), .wire_12_7_13_8_remainter(Remainder_in), .wire_13_8_14_9_remainter(Remainder_out), .wire_13_07_08_curry(C_in), .wire_13_08_09_curry(C_out));
	div_cell cas_13_7 (.~wire_out_quotient_3(T_in), .divisor[7](Divisor_in), .wire_12_6_13_7_remainter(Remainder_in), .wire_13_7_14_8_remainter(Remainder_out), .wire_13_06_07_curry(C_in), .wire_13_07_08_curry(C_out));
	div_cell cas_13_6 (.~wire_out_quotient_3(T_in), .divisor[6](Divisor_in), .wire_12_5_13_6_remainter(Remainder_in), .wire_13_6_14_7_remainter(Remainder_out), .wire_13_05_06_curry(C_in), .wire_13_06_07_curry(C_out));
	div_cell cas_13_5 (.~wire_out_quotient_3(T_in), .divisor[5](Divisor_in), .wire_12_4_13_5_remainter(Remainder_in), .wire_13_5_14_6_remainter(Remainder_out), .wire_13_04_05_curry(C_in), .wire_13_05_06_curry(C_out));
	div_cell cas_13_4 (.~wire_out_quotient_3(T_in), .divisor[4](Divisor_in), .wire_12_3_13_4_remainter(Remainder_in), .wire_13_4_14_5_remainter(Remainder_out), .wire_13_03_04_curry(C_in), .wire_13_04_05_curry(C_out));
	div_cell cas_13_3 (.~wire_out_quotient_3(T_in), .divisor[3](Divisor_in), .wire_12_2_13_3_remainter(Remainder_in), .wire_13_3_14_4_remainter(Remainder_out), .wire_13_02_03_curry(C_in), .wire_13_03_04_curry(C_out));
	div_cell cas_13_2 (.~wire_out_quotient_3(T_in), .divisor[2](Divisor_in), .wire_12_1_13_2_remainter(Remainder_in), .wire_13_2_14_3_remainter(Remainder_out), .wire_13_01_02_curry(C_in), .wire_13_02_03_curry(C_out));
	div_cell cas_13_1 (.~wire_out_quotient_3(T_in), .divisor[1](Divisor_in), .wire_12_0_13_1_remainter(Remainder_in), .wire_13_1_14_2_remainter(Remainder_out), .wire_13_00_01_curry(C_in), .wire_13_01_02_curry(C_out));
	
	div_cell cas_13_0 (.~wire_out_quotient_3(T_in), .divisor[0](Divisor_in), .dividend[3](Remainder_in), .wire_13_0_14_1_remainter(Remainder_out), .~wire_out_quotient_3(C_in), .wire_13_00_01_curry(C_out));

	//16th row
	div_cell cas_13_14 (. (T_in), . (Divisor_in), . (Remainder_in), . (Remainder_out), . (C_in), . (C_out));
	div_cell cas_13_13 ();
	div_cell cas_13_12 ();
	div_cell cas_13_11 ();
	div_cell cas_13_10 ();
	div_cell cas_13_9 ();
	div_cell cas_13_8 ();
	div_cell cas_13_7 ();
	div_cell cas_13_6 ();
	div_cell cas_13_5 ();
	div_cell cas_13_4 ();
	div_cell cas_13_3 ();
	div_cell cas_13_2 ();
	div_cell cas_13_1 ();
	div_cell cas_13_0 ();

	//17th row
	div_cell cas_13_14 (. (T_in), . (Divisor_in), . (Remainder_in), . (Remainder_out), . (C_in), . (C_out));
	div_cell cas_13_13 ();
	div_cell cas_13_12 ();
	div_cell cas_13_11 ();
	div_cell cas_13_10 ();
	div_cell cas_13_9 ();
	div_cell cas_13_8 ();
	div_cell cas_13_7 ();
	div_cell cas_13_6 ();
	div_cell cas_13_5 ();
	div_cell cas_13_4 ();
	div_cell cas_13_3 ();
	div_cell cas_13_2 ();
	div_cell cas_13_1 ();
	div_cell cas_13_0 ();

endmodule // interconect_cells