module UARTBudRateGenerator(

);

endmodule // UARTBudRateGenerator