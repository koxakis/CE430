module MAC_mac_unit(
  
);

endmodule // MAC_mac_unit