module VGASystem(
  reset,
  clk,
  VGA_Red,
  VGA_Green,
  VGA_Blue,
  VGA_HSYNC,
  VGA_VSYNC
);

input reset, clk;

output 

endmodule // VGASystem