module MAC_top_level(
  
);

endmodule // MAC_top_level