module interconect_cells(
	clk,
	reset,
	divisor,
	dividend,
	mode,
	valid_input,
	valid_output,
	final_output
);

	input [31:0] dividend;
	input [15:0] divisor;

	input clk, reset;
	input valid_input;

	output valid_output;
	output [16:0] final_output;

	assign final_output = (mode) div_res : mod_res;

	assign div_res[14] = wire_out_quotient_14;
	assign div_res[13] = wire_out_quotient_13;
	assign div_res[12] = wire_out_quotient_12;
	assign div_res[11] = wire_out_quotient_11;
	assign div_res[10] = wire_out_quotient_10;
	assign div_res[9] = wire_out_quotient_9;
	assign div_res[8] = wire_out_quotient_8;
	assign div_res[7] = wire_out_quotient_7;
	assign div_res[6] = wire_out_quotient_6;
	assign div_res[5] = wire_out_quotient_5;
	assign div_res[4] = wire_out_quotient_4;
	assign div_res[3] = wire_out_quotient_3;
	assign div_res[2] = wire_out_quotient_2;
	assign div_res[1] = wire_out_quotient_1;
	assign div_res[0] = wire_out_quotient_0;

	assign mod_res[14] = wire_out_remainder_14;
	assign mod_res[13] = wire_out_remainder_13;
	assign mod_res[12] = wire_out_remainder_12;
	assign mod_res[11] = wire_out_remainder_11;
	assign mod_res[10] = wire_out_remainder_10;
	assign mod_res[9] = wire_out_remainder_9;
	assign mod_res[8] = wire_out_remainder_8;
	assign mod_res[7] = wire_out_remainder_7;
	assign mod_res[6] = wire_out_remainder_6;
	assign mod_res[5] = wire_out_remainder_5;
	assign mod_res[4] = wire_out_remainder_4;
	assign mod_res[3] = wire_out_remainder_3;
	assign mod_res[2] = wire_out_remainder_2;
	assign mod_res[1] = wire_out_remainder_1;
	assign mod_res[0] = wire_out_remainder_0;	

	//div_cell cas_X_Y (clk,reset,T_in,Divisor_in,Remainder_in/dividend,Remainder_out,C_in,C_out);
	//1st row
	div_cell cas_0_14 (.clk(clk), .reset(reset), .1'b1(T_in), .divisor[14](Divisor_in), .dividend[30](Remainder_in), .wire_out_quotient_14(Remainder_out), .wire_13_14_curry(C_in), .(C_out) );
	div_cell cas_0_13 (.clk(clk), .reset(reset), .1'b1(T_in), .divisor[13](Divisor_in), .dividend[29](Remainder_in), .wire_0_13_1_13_remainter(Remainder_out), .wire_12_13_curry(C_in), .wire_13_14_curry(C_out) );
	div_cell cas_0_12 (.clk(clk), .reset(reset), .1'b1(T_in), .divisor[12](Divisor_in), .dividend[28](Remainder_in), .wire_0_12_1_12_remainter(Remainder_out), .wire_11_12_curry(C_in), .wire_12_13_curry(C_out) );
	div_cell cas_0_11 (.clk(clk), .reset(reset), .1'b1(T_in), .divisor[11](Divisor_in), .dividend[27](Remainder_in), .wire_0_11_1_11_remainter(Remainder_out), .wire_10_11_curry(C_in), .wire_11_12_curry(C_out) );
	div_cell cas_0_10 (.clk(clk), .reset(reset), .1'b1(T_in), .divisor[10](Divisor_in), .dividend[26](Remainder_in), .wire_0_10_1_10_remainter(Remainder_out), .wire_09_10_curry(C_in), .wire_10_11_curry(C_out) );
	div_cell cas_0_9 (.clk(clk), .reset(reset), .1'b1(T_in), .divisor[9](Divisor_in), .dividend[25](Remainder_in), .wire_0_9_1_9_remainter(Remainder_out), .wire_08_09_curry(C_in), .wire_09_10_curry(C_out) );
	div_cell cas_0_8 (.clk(clk), .reset(reset), .1'b1(T_in), .divisor[8](Divisor_in), .dividend[24](Remainder_in), .wire_0_8_1_8_remainter(Remainder_out), .wire_07_08_curry(C_in), .wire_08_09_curry(C_out) );
	div_cell cas_0_7 (.clk(clk), .reset(reset), .1'b1(T_in), .divisor[7](Divisor_in), .dividend[23](Remainder_in), .wire_0_7_1_7_remainter(Remainder_out), .wire_06_07_curry(C_in), .wire_07_08_curry(C_out) );
	div_cell cas_0_6 (.clk(clk), .reset(reset), .1'b1(T_in), .divisor[6](Divisor_in), .dividend[22](Remainder_in), .wire_0_6_1_6_remainter(Remainder_out), .wire_05_06_curry(C_in), .wire_06_07_curry(C_out) );
	div_cell cas_0_5 (.clk(clk), .reset(reset), .1'b1(T_in), .divisor[5](Divisor_in), .dividend[21](Remainder_in), .wire_0_5_1_5_remainter(Remainder_out), .wire_04_05_curry(C_in), .wire_05_06_curry(C_out) );
	div_cell cas_0_4 (.clk(clk), .reset(reset), .1'b1(T_in), .divisor[4](Divisor_in), .dividend[20](Remainder_in), .wire_0_4_1_4_remainter(Remainder_out), .wire_03_04_curry(C_in), .wire_04_05_curry(C_out) );
	div_cell cas_0_3 (.clk(clk), .reset(reset), .1'b1(T_in), .divisor[3](Divisor_in), .dividend[19](Remainder_in), .wire_0_3_1_3_remainter(Remainder_out), .wire_02_03_curry(C_in), .wire_03_04_curry(C_out) );
	div_cell cas_0_2 (.clk(clk), .reset(reset), .1'b1(T_in), .divisor[2](Divisor_in), .dividend[18](Remainder_in), .wire_0_2_1_2_remainter(Remainder_out), .wire_01_02_curry(C_in), .wire_02_03_curry(C_out) );
	div_cell cas_0_1 (.clk(clk), .reset(reset), .1'b1(T_in), .divisor[1](Divisor_in), .dividend[17](Remainder_in), .wire_0_1_1_1_remainter(Remainder_out), .wire_00_01_curry(C_in), .wire_01_02_curry(C_out) );
	div_cell cas_0_0 (.clk(clk), .reset(reset), .1'b1(T_in), .divisor[0](Divisor_in), .dividend[16](Remainder_in), .wire_0_0_1_0_remainter(Remainder_out), .1'b1(C_in), .wire_00_01_curry(C_out) );

	//2nd row
	div_cell cas_1_13 ();
	div_cell cas_1_12 ();
	div_cell cas_1_11 ();
	div_cell cas_1_10 ();
	div_cell cas_1_9 ();
	div_cell cas_1_8 ();
	div_cell cas_1_7 ();
	div_cell cas_1_6 ();
	div_cell cas_1_5 ();
	div_cell cas_1_4 ();
	div_cell cas_1_3 ();
	div_cell cas_1_2 ();
	div_cell cas_1_1 ();
	div_cell cas_1_0 ();

	//3rd row
	div_cell cas_2_13 ();
	div_cell cas_2_12 ();
	div_cell cas_2_11 ();
	div_cell cas_2_10 ();
	div_cell cas_2_9 ();
	div_cell cas_2_8 ();
	div_cell cas_2_7 ();
	div_cell cas_2_6 ();
	div_cell cas_2_5 ();
	div_cell cas_2_4 ();
	div_cell cas_2_3 ();
	div_cell cas_2_2 ();
	div_cell cas_2_1 ();
	div_cell cas_2_0 ();

	//4th row
	div_cell cas_3_13 ();
	div_cell cas_3_12 ();
	div_cell cas_3_11 ();
	div_cell cas_3_10 ();
	div_cell cas_3_9 ();
	div_cell cas_3_8 ();
	div_cell cas_3_7 ();
	div_cell cas_3_6 ();
	div_cell cas_3_5 ();
	div_cell cas_3_4 ();
	div_cell cas_3_3 ();
	div_cell cas_3_2 ();
	div_cell cas_3_1 ();
	div_cell cas_3_0 ();

	//5th row
	div_cell cas_4_13 ();
	div_cell cas_4_12 ();
	div_cell cas_4_11 ();
	div_cell cas_4_10 ();
	div_cell cas_4_9 ();
	div_cell cas_4_8 ();
	div_cell cas_4_7 ();
	div_cell cas_4_6 ();
	div_cell cas_4_5 ();
	div_cell cas_4_4 ();
	div_cell cas_4_3 ();
	div_cell cas_4_2 ();
	div_cell cas_4_1 ();
	div_cell cas_4_0 ();

	//6th row
	div_cell cas_5_13 ();
	div_cell cas_5_12 ();
	div_cell cas_5_11 ();
	div_cell cas_5_10 ();
	div_cell cas_5_9 ();
	div_cell cas_5_8 ();
	div_cell cas_5_7 ();
	div_cell cas_5_6 ();
	div_cell cas_5_5 ();
	div_cell cas_5_4 ();
	div_cell cas_5_3 ();
	div_cell cas_5_2 ();
	div_cell cas_5_1 ();
	div_cell cas_5_0 ();

	//7th row
	div_cell cas_6_13 ();
	div_cell cas_6_12 ();
	div_cell cas_6_11 ();
	div_cell cas_6_10 ();
	div_cell cas_6_9 ();
	div_cell cas_6_8 ();
	div_cell cas_6_7 ();
	div_cell cas_6_6 ();
	div_cell cas_6_5 ();
	div_cell cas_6_4 ();
	div_cell cas_6_3 ();
	div_cell cas_6_2 ();
	div_cell cas_6_1 ();
	div_cell cas_6_0 ();

	//8th row
	div_cell cas_7_13 ();
	div_cell cas_7_12 ();
	div_cell cas_7_11 ();
	div_cell cas_7_10 ();
	div_cell cas_7_9 ();
	div_cell cas_7_8 ();
	div_cell cas_7_7 ();
	div_cell cas_7_6 ();
	div_cell cas_7_5 ();
	div_cell cas_7_4 ();
	div_cell cas_7_3 ();
	div_cell cas_7_2 ();
	div_cell cas_7_1 ();
	div_cell cas_7_0 ();

	//9th row
	div_cell cas_8_13 ();
	div_cell cas_8_12 ();
	div_cell cas_8_11 ();
	div_cell cas_8_10 ();
	div_cell cas_8_9 ();
	div_cell cas_8_8 ();
	div_cell cas_8_7 ();
	div_cell cas_8_6 ();
	div_cell cas_8_5 ();
	div_cell cas_8_4 ();
	div_cell cas_8_3 ();
	div_cell cas_8_2 ();
	div_cell cas_8_1 ();
	div_cell cas_8_0 ();

	//10th row
	div_cell cas_9_13 ();
	div_cell cas_9_12 ();
	div_cell cas_9_11 ();
	div_cell cas_9_10 ();
	div_cell cas_9_9 ();
	div_cell cas_9_8 ();
	div_cell cas_9_7 ();
	div_cell cas_9_6 ();
	div_cell cas_9_5 ();
	div_cell cas_9_4 ();
	div_cell cas_9_3 ();
	div_cell cas_9_2 ();
	div_cell cas_9_1 ();
	div_cell cas_9_0 ();

	//11th row
	div_cell cas_10_13 ();
	div_cell cas_10_12 ();
	div_cell cas_10_11 ();
	div_cell cas_10_10 ();
	div_cell cas_10_9 ();
	div_cell cas_10_8 ();
	div_cell cas_10_7 ();
	div_cell cas_10_6 ();
	div_cell cas_10_5 ();
	div_cell cas_10_4 ();
	div_cell cas_10_3 ();
	div_cell cas_10_2 ();
	div_cell cas_10_1 ();
	div_cell cas_10_0 ();

	//12th row
	div_cell cas_11_13 ();
	div_cell cas_11_12 ();
	div_cell cas_11_11 ();
	div_cell cas_11_10 ();
	div_cell cas_11_9 ();
	div_cell cas_11_8 ();
	div_cell cas_11_7 ();
	div_cell cas_11_6 ();
	div_cell cas_11_5 ();
	div_cell cas_11_4 ();
	div_cell cas_11_3 ();
	div_cell cas_11_2 ();
	div_cell cas_11_1 ();
	div_cell cas_11_0 ();

	//13th row
	div_cell cas_12_13 ();
	div_cell cas_12_12 ();
	div_cell cas_12_11 ();
	div_cell cas_12_10 ();
	div_cell cas_12_9 ();
	div_cell cas_12_8 ();
	div_cell cas_12_7 ();
	div_cell cas_12_6 ();
	div_cell cas_12_5 ();
	div_cell cas_12_4 ();
	div_cell cas_12_3 ();
	div_cell cas_12_2 ();
	div_cell cas_12_1 ();
	div_cell cas_12_0 ();

	//14th row
	div_cell cas_13_13 ();
	div_cell cas_13_12 ();
	div_cell cas_13_11 ();
	div_cell cas_13_10 ();
	div_cell cas_13_9 ();
	div_cell cas_13_8 ();
	div_cell cas_13_7 ();
	div_cell cas_13_6 ();
	div_cell cas_13_5 ();
	div_cell cas_13_4 ();
	div_cell cas_13_3 ();
	div_cell cas_13_2 ();
	div_cell cas_13_1 ();
	div_cell cas_13_0 ();

endmodule // interconect_cells