module MAC_control_unit(
  
);

endmodule // MAC_control_unit