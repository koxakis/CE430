module LEDdebouncer(
	reset,
	clk,
	rb_noise,
	rb_clean
);

endmodule // LEDdebouncer