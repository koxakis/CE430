module curry_lookahead_cell(
	clk,
	reset,

);

	

endmodule // curry_lookahead_cel	clk,
